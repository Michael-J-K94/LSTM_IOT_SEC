`timescale 1ns/100ps
`define INIT_DELAY 10
`define INTERVAL 1
`define MEM_SIZE 65536

module br_weight_memory(
	input readM,
	output reg ready,
	output reg [7:0] data
	);

	reg [7:0] memory [`MEM_SIZE - 1:0];
	reg [15:0] address;

	always begin
		#`INIT_DELAY
		forever begin
			wait(readM == 1);
			#`INTERVAL;
			data = memory[address];
			address = address + 1;
			ready = 1;
			wait(readM == 0);
			#`INTERVAL;
			ready = 0;
		end
	end

	initial begin
		address <= 0;
		ready <= 0;
	end

	initial begin
		memory[16'h0] <= 8'h67;
		memory[16'h1] <= 8'hc6;
		memory[16'h2] <= 8'h69;
		memory[16'h3] <= 8'h73;
		memory[16'h4] <= 8'h51;
		memory[16'h5] <= 8'hff;
		memory[16'h6] <= 8'h4a;
		memory[16'h7] <= 8'hec;
		memory[16'h8] <= 8'h29;
		memory[16'h9] <= 8'hcd;
		memory[16'ha] <= 8'hba;
		memory[16'hb] <= 8'hab;
		memory[16'hc] <= 8'hf2;
		memory[16'hd] <= 8'hfb;
		memory[16'he] <= 8'he3;
		memory[16'hf] <= 8'h46;
		memory[16'h10] <= 8'h7c;
		memory[16'h11] <= 8'hc2;
		memory[16'h12] <= 8'h54;
		memory[16'h13] <= 8'hf8;
		memory[16'h14] <= 8'h1b;
		memory[16'h15] <= 8'he8;
		memory[16'h16] <= 8'he7;
		memory[16'h17] <= 8'h8d;
		memory[16'h18] <= 8'h76;
		memory[16'h19] <= 8'h5a;
		memory[16'h1a] <= 8'h2e;
		memory[16'h1b] <= 8'h63;
		memory[16'h1c] <= 8'h33;
		memory[16'h1d] <= 8'h9f;
		memory[16'h1e] <= 8'hc9;
		memory[16'h1f] <= 8'h9a;
		memory[16'h20] <= 8'h66;
		memory[16'h21] <= 8'h32;
		memory[16'h22] <= 8'hd;
		memory[16'h23] <= 8'hb7;
		memory[16'h24] <= 8'h31;
		memory[16'h25] <= 8'h58;
		memory[16'h26] <= 8'ha3;
		memory[16'h27] <= 8'h5a;
		memory[16'h28] <= 8'h25;
		memory[16'h29] <= 8'h5d;
		memory[16'h2a] <= 8'h5;
		memory[16'h2b] <= 8'h17;
		memory[16'h2c] <= 8'h58;
		memory[16'h2d] <= 8'he9;
		memory[16'h2e] <= 8'h5e;
		memory[16'h2f] <= 8'hd4;
		memory[16'h30] <= 8'hab;
		memory[16'h31] <= 8'hb2;
		memory[16'h32] <= 8'hcd;
		memory[16'h33] <= 8'hc6;
		memory[16'h34] <= 8'h9b;
		memory[16'h35] <= 8'hb4;
		memory[16'h36] <= 8'h54;
		memory[16'h37] <= 8'h11;
		memory[16'h38] <= 8'he;
		memory[16'h39] <= 8'h82;
		memory[16'h3a] <= 8'h74;
		memory[16'h3b] <= 8'h41;
		memory[16'h3c] <= 8'h21;
		memory[16'h3d] <= 8'h3d;
		memory[16'h3e] <= 8'hdc;
		memory[16'h3f] <= 8'h87;
		memory[16'h40] <= 8'h70;
		memory[16'h41] <= 8'he9;
		memory[16'h42] <= 8'h3e;
		memory[16'h43] <= 8'ha1;
		memory[16'h44] <= 8'h41;
		memory[16'h45] <= 8'he1;
		memory[16'h46] <= 8'hfc;
		memory[16'h47] <= 8'h67;
		memory[16'h48] <= 8'h3e;
		memory[16'h49] <= 8'h1;
		memory[16'h4a] <= 8'h7e;
		memory[16'h4b] <= 8'h97;
		memory[16'h4c] <= 8'hea;
		memory[16'h4d] <= 8'hdc;
		memory[16'h4e] <= 8'h6b;
		memory[16'h4f] <= 8'h96;
		memory[16'h50] <= 8'h8f;
		memory[16'h51] <= 8'h38;
		memory[16'h52] <= 8'h5c;
		memory[16'h53] <= 8'h2a;
		memory[16'h54] <= 8'hec;
		memory[16'h55] <= 8'hb0;
		memory[16'h56] <= 8'h3b;
		memory[16'h57] <= 8'hfb;
		memory[16'h58] <= 8'h32;
		memory[16'h59] <= 8'haf;
		memory[16'h5a] <= 8'h3c;
		memory[16'h5b] <= 8'h54;
		memory[16'h5c] <= 8'hec;
		memory[16'h5d] <= 8'h18;
		memory[16'h5e] <= 8'hdb;
		memory[16'h5f] <= 8'h5c;
		memory[16'h60] <= 8'h2;
		memory[16'h61] <= 8'h1a;
		memory[16'h62] <= 8'hfe;
		memory[16'h63] <= 8'h43;
		memory[16'h64] <= 8'hfb;
		memory[16'h65] <= 8'hfa;
		memory[16'h66] <= 8'haa;
		memory[16'h67] <= 8'h3a;
		memory[16'h68] <= 8'hfb;
		memory[16'h69] <= 8'h29;
		memory[16'h6a] <= 8'hd1;
		memory[16'h6b] <= 8'he6;
		memory[16'h6c] <= 8'h5;
		memory[16'h6d] <= 8'h3c;
		memory[16'h6e] <= 8'h7c;
		memory[16'h6f] <= 8'h94;
		memory[16'h70] <= 8'h75;
		memory[16'h71] <= 8'hd8;
		memory[16'h72] <= 8'hbe;
		memory[16'h73] <= 8'h61;
		memory[16'h74] <= 8'h89;
		memory[16'h75] <= 8'hf9;
		memory[16'h76] <= 8'h5c;
		memory[16'h77] <= 8'hbb;
		memory[16'h78] <= 8'ha8;
		memory[16'h79] <= 8'h99;
		memory[16'h7a] <= 8'hf;
		memory[16'h7b] <= 8'h95;
		memory[16'h7c] <= 8'hb1;
		memory[16'h7d] <= 8'heb;
		memory[16'h7e] <= 8'hf1;
		memory[16'h7f] <= 8'hb3;
		memory[16'h80] <= 8'h5;
		memory[16'h81] <= 8'hef;
		memory[16'h82] <= 8'hf7;
		memory[16'h83] <= 8'h0;
		memory[16'h84] <= 8'he9;
		memory[16'h85] <= 8'ha1;
		memory[16'h86] <= 8'h3a;
		memory[16'h87] <= 8'he5;
		memory[16'h88] <= 8'hca;
		memory[16'h89] <= 8'hb;
		memory[16'h8a] <= 8'hcb;
		memory[16'h8b] <= 8'hd0;
		memory[16'h8c] <= 8'h48;
		memory[16'h8d] <= 8'h47;
		memory[16'h8e] <= 8'h64;
		memory[16'h8f] <= 8'hbd;
		memory[16'h90] <= 8'h1f;
		memory[16'h91] <= 8'h23;
		memory[16'h92] <= 8'h1e;
		memory[16'h93] <= 8'ha8;
		memory[16'h94] <= 8'h1c;
		memory[16'h95] <= 8'h7b;
		memory[16'h96] <= 8'h64;
		memory[16'h97] <= 8'hc5;
		memory[16'h98] <= 8'h14;
		memory[16'h99] <= 8'h73;
		memory[16'h9a] <= 8'h5a;
		memory[16'h9b] <= 8'hc5;
		memory[16'h9c] <= 8'h5e;
		memory[16'h9d] <= 8'h4b;
		memory[16'h9e] <= 8'h79;
		memory[16'h9f] <= 8'h63;
		memory[16'ha0] <= 8'h3b;
		memory[16'ha1] <= 8'h70;
		memory[16'ha2] <= 8'h64;
		memory[16'ha3] <= 8'h24;
		memory[16'ha4] <= 8'h11;
		memory[16'ha5] <= 8'h9e;
		memory[16'ha6] <= 8'h9;
		memory[16'ha7] <= 8'hdc;
		memory[16'ha8] <= 8'haa;
		memory[16'ha9] <= 8'hd4;
		memory[16'haa] <= 8'hac;
		memory[16'hab] <= 8'hf2;
		memory[16'hac] <= 8'h1b;
		memory[16'had] <= 8'h10;
		memory[16'hae] <= 8'haf;
		memory[16'haf] <= 8'h3b;
		memory[16'hb0] <= 8'h33;
		memory[16'hb1] <= 8'hcd;
		memory[16'hb2] <= 8'he3;
		memory[16'hb3] <= 8'h50;
		memory[16'hb4] <= 8'h48;
		memory[16'hb5] <= 8'h47;
		memory[16'hb6] <= 8'h15;
		memory[16'hb7] <= 8'h5c;
		memory[16'hb8] <= 8'hbb;
		memory[16'hb9] <= 8'h6f;
		memory[16'hba] <= 8'h22;
		memory[16'hbb] <= 8'h19;
		memory[16'hbc] <= 8'hba;
		memory[16'hbd] <= 8'h9b;
		memory[16'hbe] <= 8'h7d;
		memory[16'hbf] <= 8'hf5;
		memory[16'hc0] <= 8'hb;
		memory[16'hc1] <= 8'he1;
		memory[16'hc2] <= 8'h1a;
		memory[16'hc3] <= 8'h1c;
		memory[16'hc4] <= 8'h7f;
		memory[16'hc5] <= 8'h23;
		memory[16'hc6] <= 8'hf8;
		memory[16'hc7] <= 8'h29;
		memory[16'hc8] <= 8'hf8;
		memory[16'hc9] <= 8'ha4;
		memory[16'hca] <= 8'h1b;
		memory[16'hcb] <= 8'h13;
		memory[16'hcc] <= 8'hb5;
		memory[16'hcd] <= 8'hca;
		memory[16'hce] <= 8'h4e;
		memory[16'hcf] <= 8'he8;
		memory[16'hd0] <= 8'h98;
		memory[16'hd1] <= 8'h32;
		memory[16'hd2] <= 8'h38;
		memory[16'hd3] <= 8'he0;
		memory[16'hd4] <= 8'h79;
		memory[16'hd5] <= 8'h4d;
		memory[16'hd6] <= 8'h3d;
		memory[16'hd7] <= 8'h34;
		memory[16'hd8] <= 8'hbc;
		memory[16'hd9] <= 8'h5f;
		memory[16'hda] <= 8'h4e;
		memory[16'hdb] <= 8'h77;
		memory[16'hdc] <= 8'hfa;
		memory[16'hdd] <= 8'hcb;
		memory[16'hde] <= 8'h6c;
		memory[16'hdf] <= 8'h5;
		memory[16'he0] <= 8'hac;
		memory[16'he1] <= 8'h86;
		memory[16'he2] <= 8'h21;
		memory[16'he3] <= 8'h2b;
		memory[16'he4] <= 8'haa;
		memory[16'he5] <= 8'h1a;
		memory[16'he6] <= 8'h55;
		memory[16'he7] <= 8'ha2;
		memory[16'he8] <= 8'hbe;
		memory[16'he9] <= 8'h70;
		memory[16'hea] <= 8'hb5;
		memory[16'heb] <= 8'h73;
		memory[16'hec] <= 8'h3b;
		memory[16'hed] <= 8'h4;
		memory[16'hee] <= 8'h5c;
		memory[16'hef] <= 8'hd3;
		memory[16'hf0] <= 8'h36;
		memory[16'hf1] <= 8'h94;
		memory[16'hf2] <= 8'hb3;
		memory[16'hf3] <= 8'haf;
		memory[16'hf4] <= 8'he2;
		memory[16'hf5] <= 8'hf0;
		memory[16'hf6] <= 8'he4;
		memory[16'hf7] <= 8'h9e;
		memory[16'hf8] <= 8'h4f;
		memory[16'hf9] <= 8'h32;
		memory[16'hfa] <= 8'h15;
		memory[16'hfb] <= 8'h49;
		memory[16'hfc] <= 8'hfd;
		memory[16'hfd] <= 8'h82;
		memory[16'hfe] <= 8'h4e;
		memory[16'hff] <= 8'ha9;
		memory[16'h100] <= 8'h8;
		memory[16'h101] <= 8'h70;
		memory[16'h102] <= 8'hd4;
		memory[16'h103] <= 8'hb2;
		memory[16'h104] <= 8'h8a;
		memory[16'h105] <= 8'h29;
		memory[16'h106] <= 8'h54;
		memory[16'h107] <= 8'h48;
		memory[16'h108] <= 8'h9a;
		memory[16'h109] <= 8'ha;
		memory[16'h10a] <= 8'hbc;
		memory[16'h10b] <= 8'hd5;
		memory[16'h10c] <= 8'he;
		memory[16'h10d] <= 8'h18;
		memory[16'h10e] <= 8'ha8;
		memory[16'h10f] <= 8'h44;
		memory[16'h110] <= 8'hac;
		memory[16'h111] <= 8'h5b;
		memory[16'h112] <= 8'hf3;
		memory[16'h113] <= 8'h8e;
		memory[16'h114] <= 8'h4c;
		memory[16'h115] <= 8'hd7;
		memory[16'h116] <= 8'h2d;
		memory[16'h117] <= 8'h9b;
		memory[16'h118] <= 8'h9;
		memory[16'h119] <= 8'h42;
		memory[16'h11a] <= 8'he5;
		memory[16'h11b] <= 8'h6;
		memory[16'h11c] <= 8'hc4;
		memory[16'h11d] <= 8'h33;
		memory[16'h11e] <= 8'haf;
		memory[16'h11f] <= 8'hcd;
		memory[16'h120] <= 8'ha3;
		memory[16'h121] <= 8'h84;
		memory[16'h122] <= 8'h7f;
		memory[16'h123] <= 8'h2d;
		memory[16'h124] <= 8'had;
		memory[16'h125] <= 8'hd4;
		memory[16'h126] <= 8'h76;
		memory[16'h127] <= 8'h47;
		memory[16'h128] <= 8'hde;
		memory[16'h129] <= 8'h32;
		memory[16'h12a] <= 8'h1c;
		memory[16'h12b] <= 8'hec;
		memory[16'h12c] <= 8'h4a;
		memory[16'h12d] <= 8'hc4;
		memory[16'h12e] <= 8'h30;
		memory[16'h12f] <= 8'hf6;
		memory[16'h130] <= 8'h20;
		memory[16'h131] <= 8'h23;
		memory[16'h132] <= 8'h85;
		memory[16'h133] <= 8'h6c;
		memory[16'h134] <= 8'hfb;
		memory[16'h135] <= 8'hb2;
		memory[16'h136] <= 8'h7;
		memory[16'h137] <= 8'h4;
		memory[16'h138] <= 8'hf4;
		memory[16'h139] <= 8'hec;
		memory[16'h13a] <= 8'hb;
		memory[16'h13b] <= 8'hb9;
		memory[16'h13c] <= 8'h20;
		memory[16'h13d] <= 8'hba;
		memory[16'h13e] <= 8'h86;
		memory[16'h13f] <= 8'hc3;
		memory[16'h140] <= 8'h3e;
		memory[16'h141] <= 8'h5;
		memory[16'h142] <= 8'hf1;
		memory[16'h143] <= 8'hec;
		memory[16'h144] <= 8'hd9;
		memory[16'h145] <= 8'h67;
		memory[16'h146] <= 8'h33;
		memory[16'h147] <= 8'hb7;
		memory[16'h148] <= 8'h99;
		memory[16'h149] <= 8'h50;
		memory[16'h14a] <= 8'ha3;
		memory[16'h14b] <= 8'he3;
		memory[16'h14c] <= 8'h14;
		memory[16'h14d] <= 8'hd3;
		memory[16'h14e] <= 8'hd9;
		memory[16'h14f] <= 8'h34;
		memory[16'h150] <= 8'hf7;
		memory[16'h151] <= 8'h5e;
		memory[16'h152] <= 8'ha0;
		memory[16'h153] <= 8'hf2;
		memory[16'h154] <= 8'h10;
		memory[16'h155] <= 8'ha8;
		memory[16'h156] <= 8'hf6;
		memory[16'h157] <= 8'h5;
		memory[16'h158] <= 8'h94;
		memory[16'h159] <= 8'h1;
		memory[16'h15a] <= 8'hbe;
		memory[16'h15b] <= 8'hb4;
		memory[16'h15c] <= 8'hbc;
		memory[16'h15d] <= 8'h44;
		memory[16'h15e] <= 8'h78;
		memory[16'h15f] <= 8'hfa;
		memory[16'h160] <= 8'h49;
		memory[16'h161] <= 8'h69;
		memory[16'h162] <= 8'he6;
		memory[16'h163] <= 8'h23;
		memory[16'h164] <= 8'hd0;
		memory[16'h165] <= 8'h1a;
		memory[16'h166] <= 8'hda;
		memory[16'h167] <= 8'h69;
		memory[16'h168] <= 8'h6a;
		memory[16'h169] <= 8'h7e;
		memory[16'h16a] <= 8'h4c;
		memory[16'h16b] <= 8'h7e;
		memory[16'h16c] <= 8'h51;
		memory[16'h16d] <= 8'h25;
		memory[16'h16e] <= 8'hb3;
		memory[16'h16f] <= 8'h48;
		memory[16'h170] <= 8'h84;
		memory[16'h171] <= 8'h53;
		memory[16'h172] <= 8'h3a;
		memory[16'h173] <= 8'h94;
		memory[16'h174] <= 8'hfb;
		memory[16'h175] <= 8'h31;
		memory[16'h176] <= 8'h99;
		memory[16'h177] <= 8'h90;
		memory[16'h178] <= 8'h32;
		memory[16'h179] <= 8'h57;
		memory[16'h17a] <= 8'h44;
		memory[16'h17b] <= 8'hee;
		memory[16'h17c] <= 8'h9b;
		memory[16'h17d] <= 8'hbc;
		memory[16'h17e] <= 8'he9;
		memory[16'h17f] <= 8'he5;
		memory[16'h180] <= 8'h25;
		memory[16'h181] <= 8'hcf;
		memory[16'h182] <= 8'h8;
		memory[16'h183] <= 8'hf5;
		memory[16'h184] <= 8'he9;
		memory[16'h185] <= 8'he2;
		memory[16'h186] <= 8'h5e;
		memory[16'h187] <= 8'h53;
		memory[16'h188] <= 8'h60;
		memory[16'h189] <= 8'haa;
		memory[16'h18a] <= 8'hd2;
		memory[16'h18b] <= 8'hb2;
		memory[16'h18c] <= 8'hd0;
		memory[16'h18d] <= 8'h85;
		memory[16'h18e] <= 8'hfa;
		memory[16'h18f] <= 8'h54;
		memory[16'h190] <= 8'hd8;
		memory[16'h191] <= 8'h35;
		memory[16'h192] <= 8'he8;
		memory[16'h193] <= 8'hd4;
		memory[16'h194] <= 8'h66;
		memory[16'h195] <= 8'h82;
		memory[16'h196] <= 8'h64;
		memory[16'h197] <= 8'h98;
		memory[16'h198] <= 8'hd9;
		memory[16'h199] <= 8'ha8;
		memory[16'h19a] <= 8'h87;
		memory[16'h19b] <= 8'h75;
		memory[16'h19c] <= 8'h65;
		memory[16'h19d] <= 8'h70;
		memory[16'h19e] <= 8'h5a;
		memory[16'h19f] <= 8'h8a;
		memory[16'h1a0] <= 8'h3f;
		memory[16'h1a1] <= 8'h62;
		memory[16'h1a2] <= 8'h80;
		memory[16'h1a3] <= 8'h29;
		memory[16'h1a4] <= 8'h44;
		memory[16'h1a5] <= 8'hde;
		memory[16'h1a6] <= 8'h7c;
		memory[16'h1a7] <= 8'ha5;
		memory[16'h1a8] <= 8'h89;
		memory[16'h1a9] <= 8'h4e;
		memory[16'h1aa] <= 8'h57;
		memory[16'h1ab] <= 8'h59;
		memory[16'h1ac] <= 8'hd3;
		memory[16'h1ad] <= 8'h51;
		memory[16'h1ae] <= 8'had;
		memory[16'h1af] <= 8'hac;
		memory[16'h1b0] <= 8'h86;
		memory[16'h1b1] <= 8'h95;
		memory[16'h1b2] <= 8'h80;
		memory[16'h1b3] <= 8'hec;
		memory[16'h1b4] <= 8'h17;
		memory[16'h1b5] <= 8'he4;
		memory[16'h1b6] <= 8'h85;
		memory[16'h1b7] <= 8'hf1;
		memory[16'h1b8] <= 8'h8c;
		memory[16'h1b9] <= 8'hc;
		memory[16'h1ba] <= 8'h66;
		memory[16'h1bb] <= 8'hf1;
		memory[16'h1bc] <= 8'h7c;
		memory[16'h1bd] <= 8'hc0;
		memory[16'h1be] <= 8'h7c;
		memory[16'h1bf] <= 8'hbb;
		memory[16'h1c0] <= 8'h22;
		memory[16'h1c1] <= 8'hfc;
		memory[16'h1c2] <= 8'he4;
		memory[16'h1c3] <= 8'h66;
		memory[16'h1c4] <= 8'hda;
		memory[16'h1c5] <= 8'h61;
		memory[16'h1c6] <= 8'hb;
		memory[16'h1c7] <= 8'h63;
		memory[16'h1c8] <= 8'haf;
		memory[16'h1c9] <= 8'h62;
		memory[16'h1ca] <= 8'hbc;
		memory[16'h1cb] <= 8'h83;
		memory[16'h1cc] <= 8'hb4;
		memory[16'h1cd] <= 8'h69;
		memory[16'h1ce] <= 8'h2f;
		memory[16'h1cf] <= 8'h3a;
		memory[16'h1d0] <= 8'hff;
		memory[16'h1d1] <= 8'haf;
		memory[16'h1d2] <= 8'h27;
		memory[16'h1d3] <= 8'h16;
		memory[16'h1d4] <= 8'h93;
		memory[16'h1d5] <= 8'hac;
		memory[16'h1d6] <= 8'h7;
		memory[16'h1d7] <= 8'h1f;
		memory[16'h1d8] <= 8'hb8;
		memory[16'h1d9] <= 8'h6d;
		memory[16'h1da] <= 8'h11;
		memory[16'h1db] <= 8'h34;
		memory[16'h1dc] <= 8'h2d;
		memory[16'h1dd] <= 8'h8d;
		memory[16'h1de] <= 8'hef;
		memory[16'h1df] <= 8'h4f;
		memory[16'h1e0] <= 8'h89;
		memory[16'h1e1] <= 8'hd4;
		memory[16'h1e2] <= 8'hb6;
		memory[16'h1e3] <= 8'h63;
		memory[16'h1e4] <= 8'h35;
		memory[16'h1e5] <= 8'hc1;
		memory[16'h1e6] <= 8'hc7;
		memory[16'h1e7] <= 8'he4;
		memory[16'h1e8] <= 8'h24;
		memory[16'h1e9] <= 8'h83;
		memory[16'h1ea] <= 8'h67;
		memory[16'h1eb] <= 8'hd8;
		memory[16'h1ec] <= 8'hed;
		memory[16'h1ed] <= 8'h96;
		memory[16'h1ee] <= 8'h12;
		memory[16'h1ef] <= 8'hec;
		memory[16'h1f0] <= 8'h45;
		memory[16'h1f1] <= 8'h39;
		memory[16'h1f2] <= 8'h2;
		memory[16'h1f3] <= 8'hd8;
		memory[16'h1f4] <= 8'he5;
		memory[16'h1f5] <= 8'ha;
		memory[16'h1f6] <= 8'hf8;
		memory[16'h1f7] <= 8'h9d;
		memory[16'h1f8] <= 8'h77;
		memory[16'h1f9] <= 8'h9;
		memory[16'h1fa] <= 8'hd1;
		memory[16'h1fb] <= 8'ha5;
		memory[16'h1fc] <= 8'h96;
		memory[16'h1fd] <= 8'hc1;
		memory[16'h1fe] <= 8'hf4;
		memory[16'h1ff] <= 8'h1f;
		memory[16'h200] <= 8'h95;
		memory[16'h201] <= 8'haa;
		memory[16'h202] <= 8'h82;
		memory[16'h203] <= 8'hca;
		memory[16'h204] <= 8'h6c;
		memory[16'h205] <= 8'h49;
		memory[16'h206] <= 8'hae;
		memory[16'h207] <= 8'h90;
		memory[16'h208] <= 8'hcd;
		memory[16'h209] <= 8'h16;
		memory[16'h20a] <= 8'h68;
		memory[16'h20b] <= 8'hba;
		memory[16'h20c] <= 8'hac;
		memory[16'h20d] <= 8'h7a;
		memory[16'h20e] <= 8'ha6;
		memory[16'h20f] <= 8'hf2;
		memory[16'h210] <= 8'hb4;
		memory[16'h211] <= 8'ha8;
		memory[16'h212] <= 8'hca;
		memory[16'h213] <= 8'h99;
		memory[16'h214] <= 8'hb2;
		memory[16'h215] <= 8'hc2;
		memory[16'h216] <= 8'h37;
		memory[16'h217] <= 8'h2a;
		memory[16'h218] <= 8'hcb;
		memory[16'h219] <= 8'h8;
		memory[16'h21a] <= 8'hcf;
		memory[16'h21b] <= 8'h61;
		memory[16'h21c] <= 8'hc9;
		memory[16'h21d] <= 8'hc3;
		memory[16'h21e] <= 8'h80;
		memory[16'h21f] <= 8'h5e;
		memory[16'h220] <= 8'h6e;
		memory[16'h221] <= 8'h3;
		memory[16'h222] <= 8'h28;
		memory[16'h223] <= 8'hda;
		memory[16'h224] <= 8'h4c;
		memory[16'h225] <= 8'hd7;
		memory[16'h226] <= 8'h6a;
		memory[16'h227] <= 8'h19;
		memory[16'h228] <= 8'hed;
		memory[16'h229] <= 8'hd2;
		memory[16'h22a] <= 8'hd3;
		memory[16'h22b] <= 8'h99;
		memory[16'h22c] <= 8'h4c;
		memory[16'h22d] <= 8'h79;
		memory[16'h22e] <= 8'h8b;
		memory[16'h22f] <= 8'h0;
		memory[16'h230] <= 8'h22;
		memory[16'h231] <= 8'h56;
		memory[16'h232] <= 8'h9a;
		memory[16'h233] <= 8'hd4;
		memory[16'h234] <= 8'h18;
		memory[16'h235] <= 8'hd1;
		memory[16'h236] <= 8'hfe;
		memory[16'h237] <= 8'he4;
		memory[16'h238] <= 8'hd9;
		memory[16'h239] <= 8'hcd;
		memory[16'h23a] <= 8'h45;
		memory[16'h23b] <= 8'ha3;
		memory[16'h23c] <= 8'h91;
		memory[16'h23d] <= 8'hc6;
		memory[16'h23e] <= 8'h1;
		memory[16'h23f] <= 8'hff;
		memory[16'h240] <= 8'hc9;
		memory[16'h241] <= 8'h2a;
		memory[16'h242] <= 8'hd9;
		memory[16'h243] <= 8'h15;
		memory[16'h244] <= 8'h1;
		memory[16'h245] <= 8'h43;
		memory[16'h246] <= 8'h2f;
		memory[16'h247] <= 8'hee;
		memory[16'h248] <= 8'h15;
		memory[16'h249] <= 8'h2;
		memory[16'h24a] <= 8'h87;
		memory[16'h24b] <= 8'h61;
		memory[16'h24c] <= 8'h7c;
		memory[16'h24d] <= 8'h13;
		memory[16'h24e] <= 8'h62;
		memory[16'h24f] <= 8'h9e;
		memory[16'h250] <= 8'h69;
		memory[16'h251] <= 8'hfc;
		memory[16'h252] <= 8'h72;
		memory[16'h253] <= 8'h81;
		memory[16'h254] <= 8'hcd;
		memory[16'h255] <= 8'h71;
		memory[16'h256] <= 8'h65;
		memory[16'h257] <= 8'ha6;
		memory[16'h258] <= 8'h3e;
		memory[16'h259] <= 8'hab;
		memory[16'h25a] <= 8'h49;
		memory[16'h25b] <= 8'hcf;
		memory[16'h25c] <= 8'h71;
		memory[16'h25d] <= 8'h4b;
		memory[16'h25e] <= 8'hce;
		memory[16'h25f] <= 8'h3a;
		memory[16'h260] <= 8'h75;
		memory[16'h261] <= 8'ha7;
		memory[16'h262] <= 8'h4f;
		memory[16'h263] <= 8'h76;
		memory[16'h264] <= 8'hea;
		memory[16'h265] <= 8'h7e;
		memory[16'h266] <= 8'h64;
		memory[16'h267] <= 8'hff;
		memory[16'h268] <= 8'h81;
		memory[16'h269] <= 8'heb;
		memory[16'h26a] <= 8'h61;
		memory[16'h26b] <= 8'hfd;
		memory[16'h26c] <= 8'hfe;
		memory[16'h26d] <= 8'hc3;
		memory[16'h26e] <= 8'h9b;
		memory[16'h26f] <= 8'h67;
		memory[16'h270] <= 8'hbf;
		memory[16'h271] <= 8'hd;
		memory[16'h272] <= 8'he9;
		memory[16'h273] <= 8'h8c;
		memory[16'h274] <= 8'h7e;
		memory[16'h275] <= 8'h4e;
		memory[16'h276] <= 8'h32;
		memory[16'h277] <= 8'hbd;
		memory[16'h278] <= 8'hf9;
		memory[16'h279] <= 8'h7c;
		memory[16'h27a] <= 8'h8c;
		memory[16'h27b] <= 8'h6a;
		memory[16'h27c] <= 8'hc7;
		memory[16'h27d] <= 8'h5b;
		memory[16'h27e] <= 8'ha4;
		memory[16'h27f] <= 8'h3c;
		memory[16'h280] <= 8'h2;
		memory[16'h281] <= 8'hf4;
		memory[16'h282] <= 8'hb2;
		memory[16'h283] <= 8'hed;
		memory[16'h284] <= 8'h72;
		memory[16'h285] <= 8'h16;
		memory[16'h286] <= 8'hec;
		memory[16'h287] <= 8'hf3;
		memory[16'h288] <= 8'h1;
		memory[16'h289] <= 8'h4d;
		memory[16'h28a] <= 8'hf0;
		memory[16'h28b] <= 8'h0;
		memory[16'h28c] <= 8'h10;
		memory[16'h28d] <= 8'h8b;
		memory[16'h28e] <= 8'h67;
		memory[16'h28f] <= 8'hcf;
		memory[16'h290] <= 8'h99;
		memory[16'h291] <= 8'h50;
		memory[16'h292] <= 8'h5b;
		memory[16'h293] <= 8'h17;
		memory[16'h294] <= 8'h9f;
		memory[16'h295] <= 8'h8e;
		memory[16'h296] <= 8'hd4;
		memory[16'h297] <= 8'h98;
		memory[16'h298] <= 8'ha;
		memory[16'h299] <= 8'h61;
		memory[16'h29a] <= 8'h3;
		memory[16'h29b] <= 8'hd1;
		memory[16'h29c] <= 8'hbc;
		memory[16'h29d] <= 8'ha7;
		memory[16'h29e] <= 8'hd;
		memory[16'h29f] <= 8'hbe;
		memory[16'h2a0] <= 8'h9b;
		memory[16'h2a1] <= 8'hbf;
		memory[16'h2a2] <= 8'hab;
		memory[16'h2a3] <= 8'he;
		memory[16'h2a4] <= 8'hd5;
		memory[16'h2a5] <= 8'h98;
		memory[16'h2a6] <= 8'h1;
		memory[16'h2a7] <= 8'hd6;
		memory[16'h2a8] <= 8'he5;
		memory[16'h2a9] <= 8'hf2;
		memory[16'h2aa] <= 8'hd6;
		memory[16'h2ab] <= 8'hf6;
		memory[16'h2ac] <= 8'h7d;
		memory[16'h2ad] <= 8'h3e;
		memory[16'h2ae] <= 8'hc5;
		memory[16'h2af] <= 8'h16;
		memory[16'h2b0] <= 8'h8e;
		memory[16'h2b1] <= 8'h21;
		memory[16'h2b2] <= 8'h2e;
		memory[16'h2b3] <= 8'h2d;
		memory[16'h2b4] <= 8'haf;
		memory[16'h2b5] <= 8'h2;
		memory[16'h2b6] <= 8'hc6;
		memory[16'h2b7] <= 8'hb9;
		memory[16'h2b8] <= 8'h63;
		memory[16'h2b9] <= 8'hc9;
		memory[16'h2ba] <= 8'h8a;
		memory[16'h2bb] <= 8'h1f;
		memory[16'h2bc] <= 8'h70;
		memory[16'h2bd] <= 8'h97;
		memory[16'h2be] <= 8'hde;
		memory[16'h2bf] <= 8'hc;
		memory[16'h2c0] <= 8'h56;
		memory[16'h2c1] <= 8'h89;
		memory[16'h2c2] <= 8'h1a;
		memory[16'h2c3] <= 8'h2b;
		memory[16'h2c4] <= 8'h21;
		memory[16'h2c5] <= 8'h1b;
		memory[16'h2c6] <= 8'h1;
		memory[16'h2c7] <= 8'h7;
		memory[16'h2c8] <= 8'hd;
		memory[16'h2c9] <= 8'hd8;
		memory[16'h2ca] <= 8'hfd;
		memory[16'h2cb] <= 8'h8b;
		memory[16'h2cc] <= 8'h16;
		memory[16'h2cd] <= 8'hc2;
		memory[16'h2ce] <= 8'ha1;
		memory[16'h2cf] <= 8'ha4;
		memory[16'h2d0] <= 8'he3;
		memory[16'h2d1] <= 8'hcf;
		memory[16'h2d2] <= 8'hd2;
		memory[16'h2d3] <= 8'h92;
		memory[16'h2d4] <= 8'hd2;
		memory[16'h2d5] <= 8'h98;
		memory[16'h2d6] <= 8'h4b;
		memory[16'h2d7] <= 8'h35;
		memory[16'h2d8] <= 8'h61;
		memory[16'h2d9] <= 8'hd5;
		memory[16'h2da] <= 8'h55;
		memory[16'h2db] <= 8'hd1;
		memory[16'h2dc] <= 8'h6c;
		memory[16'h2dd] <= 8'h33;
		memory[16'h2de] <= 8'hdd;
		memory[16'h2df] <= 8'hc2;
		memory[16'h2e0] <= 8'hbc;
		memory[16'h2e1] <= 8'hf7;
		memory[16'h2e2] <= 8'hed;
		memory[16'h2e3] <= 8'hde;
		memory[16'h2e4] <= 8'h13;
		memory[16'h2e5] <= 8'hef;
		memory[16'h2e6] <= 8'he5;
		memory[16'h2e7] <= 8'h20;
		memory[16'h2e8] <= 8'hc7;
		memory[16'h2e9] <= 8'he2;
		memory[16'h2ea] <= 8'hab;
		memory[16'h2eb] <= 8'hdd;
		memory[16'h2ec] <= 8'ha4;
		memory[16'h2ed] <= 8'h4d;
		memory[16'h2ee] <= 8'h81;
		memory[16'h2ef] <= 8'h88;
		memory[16'h2f0] <= 8'h1c;
		memory[16'h2f1] <= 8'h53;
		memory[16'h2f2] <= 8'h1a;
		memory[16'h2f3] <= 8'hee;
		memory[16'h2f4] <= 8'heb;
		memory[16'h2f5] <= 8'h66;
		memory[16'h2f6] <= 8'h24;
		memory[16'h2f7] <= 8'h4c;
		memory[16'h2f8] <= 8'h3b;
		memory[16'h2f9] <= 8'h79;
		memory[16'h2fa] <= 8'h1e;
		memory[16'h2fb] <= 8'ha8;
		memory[16'h2fc] <= 8'hac;
		memory[16'h2fd] <= 8'hfb;
		memory[16'h2fe] <= 8'h6a;
		memory[16'h2ff] <= 8'h68;
		memory[16'h300] <= 8'hf3;
		memory[16'h301] <= 8'h58;
		memory[16'h302] <= 8'h46;
		memory[16'h303] <= 8'h6;
		memory[16'h304] <= 8'h47;
		memory[16'h305] <= 8'h2b;
		memory[16'h306] <= 8'h26;
		memory[16'h307] <= 8'he;
		memory[16'h308] <= 8'hd;
		memory[16'h309] <= 8'hd2;
		memory[16'h30a] <= 8'heb;
		memory[16'h30b] <= 8'hb2;
		memory[16'h30c] <= 8'h1f;
		memory[16'h30d] <= 8'h6c;
		memory[16'h30e] <= 8'h3a;
		memory[16'h30f] <= 8'h3b;
		memory[16'h310] <= 8'hc0;
		memory[16'h311] <= 8'h54;
		memory[16'h312] <= 8'h2a;
		memory[16'h313] <= 8'hab;
		memory[16'h314] <= 8'hba;
		memory[16'h315] <= 8'h4e;
		memory[16'h316] <= 8'hf8;
		memory[16'h317] <= 8'hf6;
		memory[16'h318] <= 8'hc7;
		memory[16'h319] <= 8'h16;
		memory[16'h31a] <= 8'h9e;
		memory[16'h31b] <= 8'h73;
		memory[16'h31c] <= 8'h11;
		memory[16'h31d] <= 8'h8;
		memory[16'h31e] <= 8'hdb;
		memory[16'h31f] <= 8'h4;
		memory[16'h320] <= 8'h60;
		memory[16'h321] <= 8'h22;
		memory[16'h322] <= 8'ha;
		memory[16'h323] <= 8'ha7;
		memory[16'h324] <= 8'h4d;
		memory[16'h325] <= 8'h31;
		memory[16'h326] <= 8'hb5;
		memory[16'h327] <= 8'h5b;
		memory[16'h328] <= 8'h3;
		memory[16'h329] <= 8'ha0;
		memory[16'h32a] <= 8'hd;
		memory[16'h32b] <= 8'h22;
		memory[16'h32c] <= 8'hd;
		memory[16'h32d] <= 8'h47;
		memory[16'h32e] <= 8'h5d;
		memory[16'h32f] <= 8'hcd;
		memory[16'h330] <= 8'h9b;
		memory[16'h331] <= 8'h87;
		memory[16'h332] <= 8'h78;
		memory[16'h333] <= 8'h56;
		memory[16'h334] <= 8'hd5;
		memory[16'h335] <= 8'h70;
		memory[16'h336] <= 8'h4c;
		memory[16'h337] <= 8'h9c;
		memory[16'h338] <= 8'h86;
		memory[16'h339] <= 8'hea;
		memory[16'h33a] <= 8'hf;
		memory[16'h33b] <= 8'h98;
		memory[16'h33c] <= 8'hf2;
		memory[16'h33d] <= 8'heb;
		memory[16'h33e] <= 8'h9c;
		memory[16'h33f] <= 8'h53;
		memory[16'h340] <= 8'hd;
		memory[16'h341] <= 8'ha7;
		memory[16'h342] <= 8'hfa;
		memory[16'h343] <= 8'h5a;
		memory[16'h344] <= 8'hd8;
		memory[16'h345] <= 8'hb0;
		memory[16'h346] <= 8'hb5;
		memory[16'h347] <= 8'hdb;
		memory[16'h348] <= 8'h50;
		memory[16'h349] <= 8'hc2;
		memory[16'h34a] <= 8'hfd;
		memory[16'h34b] <= 8'h5d;
		memory[16'h34c] <= 8'h9;
		memory[16'h34d] <= 8'h5a;
		memory[16'h34e] <= 8'h2a;
		memory[16'h34f] <= 8'ha5;
		memory[16'h350] <= 8'he2;
		memory[16'h351] <= 8'ha3;
		memory[16'h352] <= 8'hfb;
		memory[16'h353] <= 8'hb7;
		memory[16'h354] <= 8'h13;
		memory[16'h355] <= 8'h47;
		memory[16'h356] <= 8'h54;
		memory[16'h357] <= 8'h9a;
		memory[16'h358] <= 8'h31;
		memory[16'h359] <= 8'h63;
		memory[16'h35a] <= 8'h32;
		memory[16'h35b] <= 8'h23;
		memory[16'h35c] <= 8'h4e;
		memory[16'h35d] <= 8'hce;
		memory[16'h35e] <= 8'h76;
		memory[16'h35f] <= 8'h5b;
		memory[16'h360] <= 8'h75;
		memory[16'h361] <= 8'h71;
		memory[16'h362] <= 8'hb6;
		memory[16'h363] <= 8'h4d;
		memory[16'h364] <= 8'h21;
		memory[16'h365] <= 8'h6b;
		memory[16'h366] <= 8'h28;
		memory[16'h367] <= 8'h71;
		memory[16'h368] <= 8'h2e;
		memory[16'h369] <= 8'h25;
		memory[16'h36a] <= 8'hcf;
		memory[16'h36b] <= 8'h37;
		memory[16'h36c] <= 8'h80;
		memory[16'h36d] <= 8'hf9;
		memory[16'h36e] <= 8'hdc;
		memory[16'h36f] <= 8'h62;
		memory[16'h370] <= 8'h9c;
		memory[16'h371] <= 8'hd7;
		memory[16'h372] <= 8'h19;
		memory[16'h373] <= 8'hb0;
		memory[16'h374] <= 8'h1e;
		memory[16'h375] <= 8'h6d;
		memory[16'h376] <= 8'h4a;
		memory[16'h377] <= 8'h4f;
		memory[16'h378] <= 8'hd1;
		memory[16'h379] <= 8'h7c;
		memory[16'h37a] <= 8'h73;
		memory[16'h37b] <= 8'h1f;
		memory[16'h37c] <= 8'h4a;
		memory[16'h37d] <= 8'he9;
		memory[16'h37e] <= 8'h7b;
		memory[16'h37f] <= 8'hc0;
		memory[16'h380] <= 8'h5a;
		memory[16'h381] <= 8'h31;
		memory[16'h382] <= 8'hd;
		memory[16'h383] <= 8'h7b;
		memory[16'h384] <= 8'h9c;
		memory[16'h385] <= 8'h36;
		memory[16'h386] <= 8'hed;
		memory[16'h387] <= 8'hca;
		memory[16'h388] <= 8'h5b;
		memory[16'h389] <= 8'hbc;
		memory[16'h38a] <= 8'h2;
		memory[16'h38b] <= 8'hdb;
		memory[16'h38c] <= 8'hb5;
		memory[16'h38d] <= 8'hde;
		memory[16'h38e] <= 8'h3d;
		memory[16'h38f] <= 8'h52;
		memory[16'h390] <= 8'hb6;
		memory[16'h391] <= 8'h57;
		memory[16'h392] <= 8'h2;
		memory[16'h393] <= 8'hd4;
		memory[16'h394] <= 8'hc4;
		memory[16'h395] <= 8'h4c;
		memory[16'h396] <= 8'h24;
		memory[16'h397] <= 8'h95;
		memory[16'h398] <= 8'hc8;
		memory[16'h399] <= 8'h97;
		memory[16'h39a] <= 8'hb5;
		memory[16'h39b] <= 8'h12;
		memory[16'h39c] <= 8'h80;
		memory[16'h39d] <= 8'h30;
		memory[16'h39e] <= 8'hd2;
		memory[16'h39f] <= 8'hdb;
		memory[16'h3a0] <= 8'h61;
		memory[16'h3a1] <= 8'he0;
		memory[16'h3a2] <= 8'h56;
		memory[16'h3a3] <= 8'hfd;
		memory[16'h3a4] <= 8'h16;
		memory[16'h3a5] <= 8'h43;
		memory[16'h3a6] <= 8'hc8;
		memory[16'h3a7] <= 8'h71;
		memory[16'h3a8] <= 8'hff;
		memory[16'h3a9] <= 8'hca;
		memory[16'h3aa] <= 8'h4d;
		memory[16'h3ab] <= 8'hb5;
		memory[16'h3ac] <= 8'ha8;
		memory[16'h3ad] <= 8'h8a;
		memory[16'h3ae] <= 8'h7;
		memory[16'h3af] <= 8'h5e;
		memory[16'h3b0] <= 8'he1;
		memory[16'h3b1] <= 8'h9;
		memory[16'h3b2] <= 8'h33;
		memory[16'h3b3] <= 8'ha6;
		memory[16'h3b4] <= 8'h55;
		memory[16'h3b5] <= 8'h57;
		memory[16'h3b6] <= 8'h3b;
		memory[16'h3b7] <= 8'h1d;
		memory[16'h3b8] <= 8'hee;
		memory[16'h3b9] <= 8'hf0;
		memory[16'h3ba] <= 8'h2f;
		memory[16'h3bb] <= 8'h6e;
		memory[16'h3bc] <= 8'h20;
		memory[16'h3bd] <= 8'h2;
		memory[16'h3be] <= 8'h49;
		memory[16'h3bf] <= 8'h81;
		memory[16'h3c0] <= 8'he2;
		memory[16'h3c1] <= 8'ha0;
		memory[16'h3c2] <= 8'h7f;
		memory[16'h3c3] <= 8'hf8;
		memory[16'h3c4] <= 8'he3;
		memory[16'h3c5] <= 8'h47;
		memory[16'h3c6] <= 8'h69;
		memory[16'h3c7] <= 8'he3;
		memory[16'h3c8] <= 8'h11;
		memory[16'h3c9] <= 8'hb6;
		memory[16'h3ca] <= 8'h98;
		memory[16'h3cb] <= 8'hb9;
		memory[16'h3cc] <= 8'h41;
		memory[16'h3cd] <= 8'h9f;
		memory[16'h3ce] <= 8'h18;
		memory[16'h3cf] <= 8'h22;
		memory[16'h3d0] <= 8'ha8;
		memory[16'h3d1] <= 8'h4b;
		memory[16'h3d2] <= 8'hc8;
		memory[16'h3d3] <= 8'hfd;
		memory[16'h3d4] <= 8'ha2;
		memory[16'h3d5] <= 8'h4;
		memory[16'h3d6] <= 8'h1a;
		memory[16'h3d7] <= 8'h90;
		memory[16'h3d8] <= 8'hf4;
		memory[16'h3d9] <= 8'h49;
		memory[16'h3da] <= 8'hfe;
		memory[16'h3db] <= 8'h15;
		memory[16'h3dc] <= 8'h4b;
		memory[16'h3dd] <= 8'h48;
		memory[16'h3de] <= 8'h96;
		memory[16'h3df] <= 8'h2d;
		memory[16'h3e0] <= 8'he8;
		memory[16'h3e1] <= 8'h15;
		memory[16'h3e2] <= 8'h25;
		memory[16'h3e3] <= 8'hcb;
		memory[16'h3e4] <= 8'h5c;
		memory[16'h3e5] <= 8'h8f;
		memory[16'h3e6] <= 8'hae;
		memory[16'h3e7] <= 8'h6d;
		memory[16'h3e8] <= 8'h45;
		memory[16'h3e9] <= 8'h46;
		memory[16'h3ea] <= 8'h27;
		memory[16'h3eb] <= 8'h86;
		memory[16'h3ec] <= 8'he5;
		memory[16'h3ed] <= 8'h3f;
		memory[16'h3ee] <= 8'ha9;
		memory[16'h3ef] <= 8'h8d;
		memory[16'h3f0] <= 8'h8a;
		memory[16'h3f1] <= 8'h71;
		memory[16'h3f2] <= 8'h8a;
		memory[16'h3f3] <= 8'h2c;
		memory[16'h3f4] <= 8'h75;
		memory[16'h3f5] <= 8'ha4;
		memory[16'h3f6] <= 8'hbc;
		memory[16'h3f7] <= 8'h6a;
		memory[16'h3f8] <= 8'hee;
		memory[16'h3f9] <= 8'hba;
		memory[16'h3fa] <= 8'h7f;
		memory[16'h3fb] <= 8'h39;
		memory[16'h3fc] <= 8'h2;
		memory[16'h3fd] <= 8'h15;
		memory[16'h3fe] <= 8'h67;
		memory[16'h3ff] <= 8'hea;
		memory[16'h400] <= 8'h2b;
		memory[16'h401] <= 8'h8c;
		memory[16'h402] <= 8'hb6;
		memory[16'h403] <= 8'h87;
		memory[16'h404] <= 8'h1b;
		memory[16'h405] <= 8'h64;
		memory[16'h406] <= 8'hf5;
		memory[16'h407] <= 8'h61;
		memory[16'h408] <= 8'hab;
		memory[16'h409] <= 8'h1c;
		memory[16'h40a] <= 8'he7;
		memory[16'h40b] <= 8'h90;
		memory[16'h40c] <= 8'h5b;
		memory[16'h40d] <= 8'h90;
		memory[16'h40e] <= 8'h1e;
		memory[16'h40f] <= 8'he5;
		memory[16'h410] <= 8'h2;
		memory[16'h411] <= 8'ha8;
		memory[16'h412] <= 8'h11;
		memory[16'h413] <= 8'h77;
		memory[16'h414] <= 8'h4d;
		memory[16'h415] <= 8'hcd;
		memory[16'h416] <= 8'he1;
		memory[16'h417] <= 8'h3b;
		memory[16'h418] <= 8'h87;
		memory[16'h419] <= 8'h60;
		memory[16'h41a] <= 8'h74;
		memory[16'h41b] <= 8'h8a;
		memory[16'h41c] <= 8'h76;
		memory[16'h41d] <= 8'hdb;
		memory[16'h41e] <= 8'h74;
		memory[16'h41f] <= 8'ha1;
		memory[16'h420] <= 8'h68;
		memory[16'h421] <= 8'h2a;
		memory[16'h422] <= 8'h28;
		memory[16'h423] <= 8'h83;
		memory[16'h424] <= 8'h8f;
		memory[16'h425] <= 8'h1d;
		memory[16'h426] <= 8'he4;
		memory[16'h427] <= 8'h3a;
		memory[16'h428] <= 8'h39;
		memory[16'h429] <= 8'hcc;
		memory[16'h42a] <= 8'hca;
		memory[16'h42b] <= 8'h94;
		memory[16'h42c] <= 8'h5c;
		memory[16'h42d] <= 8'he8;
		memory[16'h42e] <= 8'h79;
		memory[16'h42f] <= 8'h5e;
		memory[16'h430] <= 8'h91;
		memory[16'h431] <= 8'h8a;
		memory[16'h432] <= 8'hd6;
		memory[16'h433] <= 8'hde;
		memory[16'h434] <= 8'h57;
		memory[16'h435] <= 8'hb7;
		memory[16'h436] <= 8'h19;
		memory[16'h437] <= 8'hdf;
		memory[16'h438] <= 8'h18;
		memory[16'h439] <= 8'h8d;
		memory[16'h43a] <= 8'h69;
		memory[16'h43b] <= 8'h8e;
		memory[16'h43c] <= 8'h69;
		memory[16'h43d] <= 8'hdd;
		memory[16'h43e] <= 8'h2f;
		memory[16'h43f] <= 8'hd1;
		memory[16'h440] <= 8'h8;
		memory[16'h441] <= 8'h57;
		memory[16'h442] <= 8'h54;
		memory[16'h443] <= 8'h97;
		memory[16'h444] <= 8'h75;
		memory[16'h445] <= 8'h39;
		memory[16'h446] <= 8'hd1;
		memory[16'h447] <= 8'hae;
		memory[16'h448] <= 8'h5;
		memory[16'h449] <= 8'h9b;
		memory[16'h44a] <= 8'h43;
		memory[16'h44b] <= 8'h61;
		memory[16'h44c] <= 8'h84;
		memory[16'h44d] <= 8'hbc;
		memory[16'h44e] <= 8'hc0;
		memory[16'h44f] <= 8'h15;
		memory[16'h450] <= 8'h47;
		memory[16'h451] <= 8'h96;
		memory[16'h452] <= 8'hf3;
		memory[16'h453] <= 8'h9e;
		memory[16'h454] <= 8'h4d;
		memory[16'h455] <= 8'hc;
		memory[16'h456] <= 8'h7d;
		memory[16'h457] <= 8'h65;
		memory[16'h458] <= 8'h99;
		memory[16'h459] <= 8'he6;
		memory[16'h45a] <= 8'hf3;
		memory[16'h45b] <= 8'h2;
		memory[16'h45c] <= 8'hc4;
		memory[16'h45d] <= 8'h22;
		memory[16'h45e] <= 8'hd3;
		memory[16'h45f] <= 8'hcc;
		memory[16'h460] <= 8'h7a;
		memory[16'h461] <= 8'h28;
		memory[16'h462] <= 8'h63;
		memory[16'h463] <= 8'hef;
		memory[16'h464] <= 8'h61;
		memory[16'h465] <= 8'h34;
		memory[16'h466] <= 8'h9d;
		memory[16'h467] <= 8'h66;
		memory[16'h468] <= 8'hcf;
		memory[16'h469] <= 8'he0;
		memory[16'h46a] <= 8'hc7;
		memory[16'h46b] <= 8'h53;
		memory[16'h46c] <= 8'h9d;
		memory[16'h46d] <= 8'h87;
		memory[16'h46e] <= 8'h68;
		memory[16'h46f] <= 8'he4;
		memory[16'h470] <= 8'h1d;
		memory[16'h471] <= 8'h5b;
		memory[16'h472] <= 8'h82;
		memory[16'h473] <= 8'h6b;
		memory[16'h474] <= 8'h67;
		memory[16'h475] <= 8'h0;
		memory[16'h476] <= 8'hd0;
		memory[16'h477] <= 8'h1;
		memory[16'h478] <= 8'he6;
		memory[16'h479] <= 8'hc4;
		memory[16'h47a] <= 8'h3;
		memory[16'h47b] <= 8'haa;
		memory[16'h47c] <= 8'he6;
		memory[16'h47d] <= 8'hd7;
		memory[16'h47e] <= 8'h76;
		memory[16'h47f] <= 8'h60;
		memory[16'h480] <= 8'hff;
		memory[16'h481] <= 8'hd9;
		memory[16'h482] <= 8'h4f;
		memory[16'h483] <= 8'h60;
		memory[16'h484] <= 8'hd;
		memory[16'h485] <= 8'hed;
		memory[16'h486] <= 8'hc6;
		memory[16'h487] <= 8'hdd;
		memory[16'h488] <= 8'hcd;
		memory[16'h489] <= 8'h8d;
		memory[16'h48a] <= 8'h30;
		memory[16'h48b] <= 8'h6a;
		memory[16'h48c] <= 8'h15;
		memory[16'h48d] <= 8'h99;
		memory[16'h48e] <= 8'h4e;
		memory[16'h48f] <= 8'h32;
		memory[16'h490] <= 8'hf4;
		memory[16'h491] <= 8'hd1;
		memory[16'h492] <= 8'h9d;
		memory[16'h493] <= 8'h5c;
		memory[16'h494] <= 8'hd1;
		memory[16'h495] <= 8'h6e;
		memory[16'h496] <= 8'h5d;
		memory[16'h497] <= 8'hb7;
		memory[16'h498] <= 8'h32;
		memory[16'h499] <= 8'h60;
		memory[16'h49a] <= 8'h62;
		memory[16'h49b] <= 8'h18;
		memory[16'h49c] <= 8'h37;
		memory[16'h49d] <= 8'hd8;
		memory[16'h49e] <= 8'h79;
		memory[16'h49f] <= 8'h36;
		memory[16'h4a0] <= 8'hb2;
		memory[16'h4a1] <= 8'hc8;
		memory[16'h4a2] <= 8'h96;
		memory[16'h4a3] <= 8'hbf;
		memory[16'h4a4] <= 8'hb5;
		memory[16'h4a5] <= 8'h5c;
		memory[16'h4a6] <= 8'h9c;
		memory[16'h4a7] <= 8'h83;
		memory[16'h4a8] <= 8'hea;
		memory[16'h4a9] <= 8'hcd;
		memory[16'h4aa] <= 8'hed;
		memory[16'h4ab] <= 8'hff;
		memory[16'h4ac] <= 8'h66;
		memory[16'h4ad] <= 8'h3c;
		memory[16'h4ae] <= 8'h31;
		memory[16'h4af] <= 8'h5a;
		memory[16'h4b0] <= 8'hd;
		memory[16'h4b1] <= 8'hcf;
		memory[16'h4b2] <= 8'hb6;
		memory[16'h4b3] <= 8'hde;
		memory[16'h4b4] <= 8'h3d;
		memory[16'h4b5] <= 8'h13;
		memory[16'h4b6] <= 8'h95;
		memory[16'h4b7] <= 8'h6f;
		memory[16'h4b8] <= 8'h74;
		memory[16'h4b9] <= 8'hf7;
		memory[16'h4ba] <= 8'h87;
		memory[16'h4bb] <= 8'hab;
		memory[16'h4bc] <= 8'hd0;
		memory[16'h4bd] <= 8'h0;
		memory[16'h4be] <= 8'he2;
		memory[16'h4bf] <= 8'h82;
		memory[16'h4c0] <= 8'hc9;
		memory[16'h4c1] <= 8'h78;
		memory[16'h4c2] <= 8'h41;
		memory[16'h4c3] <= 8'h7e;
		memory[16'h4c4] <= 8'hd5;
		memory[16'h4c5] <= 8'hde;
		memory[16'h4c6] <= 8'h1;
		memory[16'h4c7] <= 8'hbf;
		memory[16'h4c8] <= 8'hab;
		memory[16'h4c9] <= 8'hef;
		memory[16'h4ca] <= 8'hbe;
		memory[16'h4cb] <= 8'h11;
		memory[16'h4cc] <= 8'h2b;
		memory[16'h4cd] <= 8'hef;
		memory[16'h4ce] <= 8'h6b;
		memory[16'h4cf] <= 8'h38;
		memory[16'h4d0] <= 8'hbe;
		memory[16'h4d1] <= 8'h22;
		memory[16'h4d2] <= 8'h16;
		memory[16'h4d3] <= 8'hfb;
		memory[16'h4d4] <= 8'h35;
		memory[16'h4d5] <= 8'hab;
		memory[16'h4d6] <= 8'h6a;
		memory[16'h4d7] <= 8'ha9;
		memory[16'h4d8] <= 8'ha3;
		memory[16'h4d9] <= 8'hf2;
		memory[16'h4da] <= 8'h55;
		memory[16'h4db] <= 8'h73;
		memory[16'h4dc] <= 8'hf2;
		memory[16'h4dd] <= 8'h37;
		memory[16'h4de] <= 8'hf5;
		memory[16'h4df] <= 8'hbb;
		memory[16'h4e0] <= 8'haf;
		memory[16'h4e1] <= 8'h36;
		memory[16'h4e2] <= 8'h3a;
		memory[16'h4e3] <= 8'h84;
		memory[16'h4e4] <= 8'h14;
		memory[16'h4e5] <= 8'h3b;
		memory[16'h4e6] <= 8'h43;
		memory[16'h4e7] <= 8'hbf;
		memory[16'h4e8] <= 8'h2a;
		memory[16'h4e9] <= 8'h1;
		memory[16'h4ea] <= 8'hd0;
		memory[16'h4eb] <= 8'h55;
		memory[16'h4ec] <= 8'hf1;
		memory[16'h4ed] <= 8'h3c;
		memory[16'h4ee] <= 8'h8d;
		memory[16'h4ef] <= 8'haf;
		memory[16'h4f0] <= 8'h5e;
		memory[16'h4f1] <= 8'ha3;
		memory[16'h4f2] <= 8'hab;
		memory[16'h4f3] <= 8'h93;
		memory[16'h4f4] <= 8'h4f;
		memory[16'h4f5] <= 8'h15;
		memory[16'h4f6] <= 8'h3d;
		memory[16'h4f7] <= 8'hf2;
		memory[16'h4f8] <= 8'h7;
		memory[16'h4f9] <= 8'h92;
		memory[16'h4fa] <= 8'h65;
		memory[16'h4fb] <= 8'hfa;
		memory[16'h4fc] <= 8'hc9;
		memory[16'h4fd] <= 8'h5a;
		memory[16'h4fe] <= 8'hb5;
		memory[16'h4ff] <= 8'h78;
		memory[16'h500] <= 8'h90;
		memory[16'h501] <= 8'hef;
		memory[16'h502] <= 8'hfd;
		memory[16'h503] <= 8'ha5;
		memory[16'h504] <= 8'h2b;
		memory[16'h505] <= 8'h40;
		memory[16'h506] <= 8'h64;
		memory[16'h507] <= 8'h55;
		memory[16'h508] <= 8'h42;
		memory[16'h509] <= 8'h35;
		memory[16'h50a] <= 8'hab;
		memory[16'h50b] <= 8'h33;
		memory[16'h50c] <= 8'h71;
		memory[16'h50d] <= 8'h38;
		memory[16'h50e] <= 8'he2;
		memory[16'h50f] <= 8'hcf;
		memory[16'h510] <= 8'hdc;
		memory[16'h511] <= 8'h8d;
		memory[16'h512] <= 8'h62;
		memory[16'h513] <= 8'h2b;
		memory[16'h514] <= 8'ha3;
		memory[16'h515] <= 8'h9f;
		memory[16'h516] <= 8'h1d;
		memory[16'h517] <= 8'haa;
		memory[16'h518] <= 8'h31;
		memory[16'h519] <= 8'h82;
		memory[16'h51a] <= 8'ha4;
		memory[16'h51b] <= 8'hfa;
		memory[16'h51c] <= 8'hdc;
		memory[16'h51d] <= 8'h5a;
		memory[16'h51e] <= 8'h73;
		memory[16'h51f] <= 8'h6c;
		memory[16'h520] <= 8'h49;
		memory[16'h521] <= 8'h70;
		memory[16'h522] <= 8'h11;
		memory[16'h523] <= 8'h74;
		memory[16'h524] <= 8'hb0;
		memory[16'h525] <= 8'h76;
		memory[16'h526] <= 8'hca;
		memory[16'h527] <= 8'hf2;
		memory[16'h528] <= 8'hab;
		memory[16'h529] <= 8'h75;
		memory[16'h52a] <= 8'h25;
		memory[16'h52b] <= 8'h1c;
		memory[16'h52c] <= 8'had;
		memory[16'h52d] <= 8'h8;
		memory[16'h52e] <= 8'heb;
		memory[16'h52f] <= 8'h89;
		memory[16'h530] <= 8'h95;
		memory[16'h531] <= 8'h4d;
		memory[16'h532] <= 8'hb4;
		memory[16'h533] <= 8'h38;
		memory[16'h534] <= 8'hed;
		memory[16'h535] <= 8'hd1;
		memory[16'h536] <= 8'he3;
		memory[16'h537] <= 8'h1e;
		memory[16'h538] <= 8'h53;
		memory[16'h539] <= 8'h87;
		memory[16'h53a] <= 8'h19;
		memory[16'h53b] <= 8'h2f;
		memory[16'h53c] <= 8'he1;
		memory[16'h53d] <= 8'h8c;
		memory[16'h53e] <= 8'h9c;
		memory[16'h53f] <= 8'h2b;
		memory[16'h540] <= 8'hfc;
		memory[16'h541] <= 8'had;
		memory[16'h542] <= 8'h9f;
		memory[16'h543] <= 8'hac;
		memory[16'h544] <= 8'h23;
		memory[16'h545] <= 8'h69;
		memory[16'h546] <= 8'h9f;
		memory[16'h547] <= 8'hce;
		memory[16'h548] <= 8'hde;
		memory[16'h549] <= 8'hc4;
		memory[16'h54a] <= 8'hea;
		memory[16'h54b] <= 8'h8c;
		memory[16'h54c] <= 8'hcc;
		memory[16'h54d] <= 8'hd5;
		memory[16'h54e] <= 8'h15;
		memory[16'h54f] <= 8'h62;
		memory[16'h550] <= 8'h23;
		memory[16'h551] <= 8'hca;
		memory[16'h552] <= 8'h9a;
		memory[16'h553] <= 8'h10;
		memory[16'h554] <= 8'h9b;
		memory[16'h555] <= 8'h7d;
		memory[16'h556] <= 8'h2e;
		memory[16'h557] <= 8'hef;
		memory[16'h558] <= 8'h5;
		memory[16'h559] <= 8'h47;
		memory[16'h55a] <= 8'h1e;
		memory[16'h55b] <= 8'he6;
		memory[16'h55c] <= 8'hd3;
		memory[16'h55d] <= 8'hba;
		memory[16'h55e] <= 8'h11;
		memory[16'h55f] <= 8'hcf;
		memory[16'h560] <= 8'h68;
		memory[16'h561] <= 8'hb1;
		memory[16'h562] <= 8'h7c;
		memory[16'h563] <= 8'h8b;
		memory[16'h564] <= 8'h1a;
		memory[16'h565] <= 8'h1b;
		memory[16'h566] <= 8'h5a;
		memory[16'h567] <= 8'hf9;
		memory[16'h568] <= 8'hdf;
		memory[16'h569] <= 8'h44;
		memory[16'h56a] <= 8'h85;
		memory[16'h56b] <= 8'hac;
		memory[16'h56c] <= 8'h1a;
		memory[16'h56d] <= 8'h9a;
		memory[16'h56e] <= 8'he;
		memory[16'h56f] <= 8'h3d;
		memory[16'h570] <= 8'h64;
		memory[16'h571] <= 8'ha8;
		memory[16'h572] <= 8'h4d;
		memory[16'h573] <= 8'h0;
		memory[16'h574] <= 8'h26;
		memory[16'h575] <= 8'h7b;
		memory[16'h576] <= 8'hef;
		memory[16'h577] <= 8'h2b;
		memory[16'h578] <= 8'hc3;
		memory[16'h579] <= 8'hd;
		memory[16'h57a] <= 8'h11;
		memory[16'h57b] <= 8'h96;
		memory[16'h57c] <= 8'hc8;
		memory[16'h57d] <= 8'h23;
		memory[16'h57e] <= 8'h66;
		memory[16'h57f] <= 8'h30;
		memory[16'h580] <= 8'hd4;
		memory[16'h581] <= 8'he2;
		memory[16'h582] <= 8'hbb;
		memory[16'h583] <= 8'hee;
		memory[16'h584] <= 8'hfd;
		memory[16'h585] <= 8'h15;
		memory[16'h586] <= 8'he7;
		memory[16'h587] <= 8'hdc;
		memory[16'h588] <= 8'h5a;
		memory[16'h589] <= 8'h6c;
		memory[16'h58a] <= 8'h88;
		memory[16'h58b] <= 8'h74;
		memory[16'h58c] <= 8'h7;
		memory[16'h58d] <= 8'h96;
		memory[16'h58e] <= 8'hb1;
		memory[16'h58f] <= 8'h6b;
		memory[16'h590] <= 8'h3f;
		memory[16'h591] <= 8'hfe;
		memory[16'h592] <= 8'h6b;
		memory[16'h593] <= 8'h65;
		memory[16'h594] <= 8'h79;
		memory[16'h595] <= 8'h5a;
		memory[16'h596] <= 8'h90;
		memory[16'h597] <= 8'h3c;
		memory[16'h598] <= 8'h68;
		memory[16'h599] <= 8'ha1;
		memory[16'h59a] <= 8'hd3;
		memory[16'h59b] <= 8'h30;
		memory[16'h59c] <= 8'hc4;
		memory[16'h59d] <= 8'h39;
		memory[16'h59e] <= 8'h60;
		memory[16'h59f] <= 8'h98;
		memory[16'h5a0] <= 8'h1b;
		memory[16'h5a1] <= 8'h1b;
		memory[16'h5a2] <= 8'h87;
		memory[16'h5a3] <= 8'h18;
		memory[16'h5a4] <= 8'h31;
		memory[16'h5a5] <= 8'h6e;
		memory[16'h5a6] <= 8'hf4;
		memory[16'h5a7] <= 8'h8b;
		memory[16'h5a8] <= 8'hdb;
		memory[16'h5a9] <= 8'h7d;
		memory[16'h5aa] <= 8'hff;
		memory[16'h5ab] <= 8'he2;
		memory[16'h5ac] <= 8'h13;
		memory[16'h5ad] <= 8'hb0;
		memory[16'h5ae] <= 8'h4d;
		memory[16'h5af] <= 8'h52;
		memory[16'h5b0] <= 8'hae;
		memory[16'h5b1] <= 8'hb9;
		memory[16'h5b2] <= 8'hb7;
		memory[16'h5b3] <= 8'h27;
		memory[16'h5b4] <= 8'h13;
		memory[16'h5b5] <= 8'h47;
		memory[16'h5b6] <= 8'h64;
		memory[16'h5b7] <= 8'h7b;
		memory[16'h5b8] <= 8'he9;
		memory[16'h5b9] <= 8'h37;
		memory[16'h5ba] <= 8'hab;
		memory[16'h5bb] <= 8'had;
		memory[16'h5bc] <= 8'h70;
		memory[16'h5bd] <= 8'hb;
		memory[16'h5be] <= 8'h46;
		memory[16'h5bf] <= 8'h8b;
		memory[16'h5c0] <= 8'h27;
		memory[16'h5c1] <= 8'hcd;
		memory[16'h5c2] <= 8'ha3;
		memory[16'h5c3] <= 8'h58;
		memory[16'h5c4] <= 8'h3b;
		memory[16'h5c5] <= 8'h97;
		memory[16'h5c6] <= 8'he3;
		memory[16'h5c7] <= 8'h16;
		memory[16'h5c8] <= 8'h14;
		memory[16'h5c9] <= 8'he2;
		memory[16'h5ca] <= 8'hf8;
		memory[16'h5cb] <= 8'h28;
		memory[16'h5cc] <= 8'h92;
		memory[16'h5cd] <= 8'h46;
		memory[16'h5ce] <= 8'h7a;
		memory[16'h5cf] <= 8'h40;
		memory[16'h5d0] <= 8'hff;
		memory[16'h5d1] <= 8'h32;
		memory[16'h5d2] <= 8'h67;
		memory[16'h5d3] <= 8'h12;
		memory[16'h5d4] <= 8'h79;
		memory[16'h5d5] <= 8'hcb;
		memory[16'h5d6] <= 8'h8e;
		memory[16'h5d7] <= 8'h62;
		memory[16'h5d8] <= 8'h2;
		memory[16'h5d9] <= 8'h39;
		memory[16'h5da] <= 8'h10;
		memory[16'h5db] <= 8'h72;
		memory[16'h5dc] <= 8'h45;
		memory[16'h5dd] <= 8'h56;
		memory[16'h5de] <= 8'hfd;
		memory[16'h5df] <= 8'h6c;
		memory[16'h5e0] <= 8'h23;
		memory[16'h5e1] <= 8'ha0;
		memory[16'h5e2] <= 8'hc4;
		memory[16'h5e3] <= 8'h5e;
		memory[16'h5e4] <= 8'h38;
		memory[16'h5e5] <= 8'ha7;
		memory[16'h5e6] <= 8'h75;
		memory[16'h5e7] <= 8'h4c;
		memory[16'h5e8] <= 8'h89;
		memory[16'h5e9] <= 8'h6d;
		memory[16'h5ea] <= 8'h74;
		memory[16'h5eb] <= 8'h1b;
		memory[16'h5ec] <= 8'hb3;
		memory[16'h5ed] <= 8'hef;
		memory[16'h5ee] <= 8'h5b;
		memory[16'h5ef] <= 8'hb2;
		memory[16'h5f0] <= 8'h21;
		memory[16'h5f1] <= 8'hc2;
		memory[16'h5f2] <= 8'hc5;
		memory[16'h5f3] <= 8'h9a;
		memory[16'h5f4] <= 8'h8e;
		memory[16'h5f5] <= 8'h53;
		memory[16'h5f6] <= 8'hfd;
		memory[16'h5f7] <= 8'h90;
		memory[16'h5f8] <= 8'h8c;
		memory[16'h5f9] <= 8'hd;
		memory[16'h5fa] <= 8'h3;
		memory[16'h5fb] <= 8'hd1;
		memory[16'h5fc] <= 8'h63;
		memory[16'h5fd] <= 8'h0;
		memory[16'h5fe] <= 8'h3d;
		memory[16'h5ff] <= 8'h86;
		memory[16'h600] <= 8'ha1;
		memory[16'h601] <= 8'h1;
		memory[16'h602] <= 8'he4;
		memory[16'h603] <= 8'hd9;
		memory[16'h604] <= 8'ha8;
		memory[16'h605] <= 8'h59;
		memory[16'h606] <= 8'h25;
		memory[16'h607] <= 8'h31;
		memory[16'h608] <= 8'hc7;
		memory[16'h609] <= 8'h9a;
		memory[16'h60a] <= 8'h4c;
		memory[16'h60b] <= 8'h7a;
		memory[16'h60c] <= 8'h89;
		memory[16'h60d] <= 8'ha7;
		memory[16'h60e] <= 8'h2d;
		memory[16'h60f] <= 8'haa;
		memory[16'h610] <= 8'h6a;
		memory[16'h611] <= 8'hf2;
		memory[16'h612] <= 8'h44;
		memory[16'h613] <= 8'hf8;
		memory[16'h614] <= 8'h45;
		memory[16'h615] <= 8'h41;
		memory[16'h616] <= 8'h88;
		memory[16'h617] <= 8'hd1;
		memory[16'h618] <= 8'h4e;
		memory[16'h619] <= 8'h8b;
		memory[16'h61a] <= 8'ha3;
		memory[16'h61b] <= 8'hb1;
		memory[16'h61c] <= 8'h8c;
		memory[16'h61d] <= 8'he0;
		memory[16'h61e] <= 8'h37;
		memory[16'h61f] <= 8'h2d;
		memory[16'h620] <= 8'he2;
		memory[16'h621] <= 8'h1c;
		memory[16'h622] <= 8'h6;
		memory[16'h623] <= 8'h8a;
		memory[16'h624] <= 8'h75;
		memory[16'h625] <= 8'h2b;
		memory[16'h626] <= 8'hbc;
		memory[16'h627] <= 8'h3c;
		memory[16'h628] <= 8'hc5;
		memory[16'h629] <= 8'h8;
		memory[16'h62a] <= 8'hb7;
		memory[16'h62b] <= 8'h4e;
		memory[16'h62c] <= 8'hb0;
		memory[16'h62d] <= 8'he4;
		memory[16'h62e] <= 8'hf8;
		memory[16'h62f] <= 8'h1a;
		memory[16'h630] <= 8'hd6;
		memory[16'h631] <= 8'h3d;
		memory[16'h632] <= 8'h12;
		memory[16'h633] <= 8'h1b;
		memory[16'h634] <= 8'h7e;
		memory[16'h635] <= 8'h9a;
		memory[16'h636] <= 8'hec;
		memory[16'h637] <= 8'hcd;
		memory[16'h638] <= 8'h26;
		memory[16'h639] <= 8'h8f;
		memory[16'h63a] <= 8'h7e;
		memory[16'h63b] <= 8'hb2;
		memory[16'h63c] <= 8'h70;
		memory[16'h63d] <= 8'hb6;
		memory[16'h63e] <= 8'hdf;
		memory[16'h63f] <= 8'h52;
		memory[16'h640] <= 8'hd2;
		memory[16'h641] <= 8'he5;
		memory[16'h642] <= 8'hdc;
		memory[16'h643] <= 8'h47;
		memory[16'h644] <= 8'h10;
		memory[16'h645] <= 8'h98;
		memory[16'h646] <= 8'h84;
		memory[16'h647] <= 8'hd6;
		memory[16'h648] <= 8'ha1;
		memory[16'h649] <= 8'h3b;
		memory[16'h64a] <= 8'h24;
		memory[16'h64b] <= 8'h51;
		memory[16'h64c] <= 8'h1f;
		memory[16'h64d] <= 8'h1d;
		memory[16'h64e] <= 8'h6b;
		memory[16'h64f] <= 8'hf5;
		memory[16'h650] <= 8'h5a;
		memory[16'h651] <= 8'h7d;
		memory[16'h652] <= 8'h10;
		memory[16'h653] <= 8'hd8;
		memory[16'h654] <= 8'h17;
		memory[16'h655] <= 8'hfc;
		memory[16'h656] <= 8'ha5;
		memory[16'h657] <= 8'h3d;
		memory[16'h658] <= 8'h8c;
		memory[16'h659] <= 8'h24;
		memory[16'h65a] <= 8'hef;
		memory[16'h65b] <= 8'hfc;
		memory[16'h65c] <= 8'hda;
		memory[16'h65d] <= 8'hce;
		memory[16'h65e] <= 8'h4e;
		memory[16'h65f] <= 8'hac;
		memory[16'h660] <= 8'hb3;
		memory[16'h661] <= 8'h2a;
		memory[16'h662] <= 8'hf3;
		memory[16'h663] <= 8'hc4;
		memory[16'h664] <= 8'hc3;
		memory[16'h665] <= 8'h77;
		memory[16'h666] <= 8'h9a;
		memory[16'h667] <= 8'h64;
		memory[16'h668] <= 8'hb2;
		memory[16'h669] <= 8'hbe;
		memory[16'h66a] <= 8'hb5;
		memory[16'h66b] <= 8'hd1;
		memory[16'h66c] <= 8'hdb;
		memory[16'h66d] <= 8'h20;
		memory[16'h66e] <= 8'hc6;
		memory[16'h66f] <= 8'h35;
		memory[16'h670] <= 8'h9d;
		memory[16'h671] <= 8'hd6;
		memory[16'h672] <= 8'he;
		memory[16'h673] <= 8'hb4;
		memory[16'h674] <= 8'hd3;
		memory[16'h675] <= 8'hb3;
		memory[16'h676] <= 8'hf2;
		memory[16'h677] <= 8'h5f;
		memory[16'h678] <= 8'hd7;
		memory[16'h679] <= 8'he1;
		memory[16'h67a] <= 8'h5b;
		memory[16'h67b] <= 8'hb1;
		memory[16'h67c] <= 8'hb0;
		memory[16'h67d] <= 8'ha9;
		memory[16'h67e] <= 8'h5d;
		memory[16'h67f] <= 8'h63;
		memory[16'h680] <= 8'hd3;
		memory[16'h681] <= 8'h51;
		memory[16'h682] <= 8'h27;
		memory[16'h683] <= 8'h96;
		memory[16'h684] <= 8'hc8;
		memory[16'h685] <= 8'hc1;
		memory[16'h686] <= 8'hfa;
		memory[16'h687] <= 8'h7b;
		memory[16'h688] <= 8'h80;
		memory[16'h689] <= 8'haf;
		memory[16'h68a] <= 8'h4c;
		memory[16'h68b] <= 8'h5b;
		memory[16'h68c] <= 8'hcf;
		memory[16'h68d] <= 8'h13;
		memory[16'h68e] <= 8'h91;
		memory[16'h68f] <= 8'h6c;
		memory[16'h690] <= 8'he9;
		memory[16'h691] <= 8'h9f;
		memory[16'h692] <= 8'h21;
		memory[16'h693] <= 8'hbc;
		memory[16'h694] <= 8'h52;
		memory[16'h695] <= 8'h13;
		memory[16'h696] <= 8'h1b;
		memory[16'h697] <= 8'h2a;
		memory[16'h698] <= 8'hf4;
		memory[16'h699] <= 8'h76;
		memory[16'h69a] <= 8'hdb;
		memory[16'h69b] <= 8'ha4;
		memory[16'h69c] <= 8'h1f;
		memory[16'h69d] <= 8'h39;
		memory[16'h69e] <= 8'h8;
		memory[16'h69f] <= 8'hf3;
		memory[16'h6a0] <= 8'h8a;
		memory[16'h6a1] <= 8'h2f;
		memory[16'h6a2] <= 8'h89;
		memory[16'h6a3] <= 8'h52;
		memory[16'h6a4] <= 8'hf1;
		memory[16'h6a5] <= 8'h84;
		memory[16'h6a6] <= 8'hcd;
		memory[16'h6a7] <= 8'h71;
		memory[16'h6a8] <= 8'h33;
		memory[16'h6a9] <= 8'h1a;
		memory[16'h6aa] <= 8'hcc;
		memory[16'h6ab] <= 8'h3;
		memory[16'h6ac] <= 8'h2d;
		memory[16'h6ad] <= 8'h5d;
		memory[16'h6ae] <= 8'h6f;
		memory[16'h6af] <= 8'h16;
		memory[16'h6b0] <= 8'hfc;
		memory[16'h6b1] <= 8'h90;
		memory[16'h6b2] <= 8'hd3;
		memory[16'h6b3] <= 8'h4f;
		memory[16'h6b4] <= 8'ha3;
		memory[16'h6b5] <= 8'hee;
		memory[16'h6b6] <= 8'h79;
		memory[16'h6b7] <= 8'h98;
		memory[16'h6b8] <= 8'h65;
		memory[16'h6b9] <= 8'h54;
		memory[16'h6ba] <= 8'h3c;
		memory[16'h6bb] <= 8'h84;
		memory[16'h6bc] <= 8'h8d;
		memory[16'h6bd] <= 8'h44;
		memory[16'h6be] <= 8'h77;
		memory[16'h6bf] <= 8'h17;
		memory[16'h6c0] <= 8'h74;
		memory[16'h6c1] <= 8'h1;
		memory[16'h6c2] <= 8'h6a;
		memory[16'h6c3] <= 8'h65;
		memory[16'h6c4] <= 8'h85;
		memory[16'h6c5] <= 8'h37;
		memory[16'h6c6] <= 8'hd6;
		memory[16'h6c7] <= 8'hb8;
		memory[16'h6c8] <= 8'h51;
		memory[16'h6c9] <= 8'ha2;
		memory[16'h6ca] <= 8'hbb;
		memory[16'h6cb] <= 8'h7e;
		memory[16'h6cc] <= 8'h0;
		memory[16'h6cd] <= 8'h2b;
		memory[16'h6ce] <= 8'h95;
		memory[16'h6cf] <= 8'hfc;
		memory[16'h6d0] <= 8'hbb;
		memory[16'h6d1] <= 8'h68;
		memory[16'h6d2] <= 8'h4b;
		memory[16'h6d3] <= 8'h5f;
		memory[16'h6d4] <= 8'h56;
		memory[16'h6d5] <= 8'hc4;
		memory[16'h6d6] <= 8'hf7;
		memory[16'h6d7] <= 8'hbb;
		memory[16'h6d8] <= 8'h19;
		memory[16'h6d9] <= 8'h33;
		memory[16'h6da] <= 8'h40;
		memory[16'h6db] <= 8'ha6;
		memory[16'h6dc] <= 8'h78;
		memory[16'h6dd] <= 8'hb7;
		memory[16'h6de] <= 8'hbe;
		memory[16'h6df] <= 8'hec;
		memory[16'h6e0] <= 8'hb8;
		memory[16'h6e1] <= 8'h28;
		memory[16'h6e2] <= 8'h51;
		memory[16'h6e3] <= 8'h3d;
		memory[16'h6e4] <= 8'h5f;
		memory[16'h6e5] <= 8'h27;
		memory[16'h6e6] <= 8'hf6;
		memory[16'h6e7] <= 8'hb1;
		memory[16'h6e8] <= 8'hc9;
		memory[16'h6e9] <= 8'hb1;
		memory[16'h6ea] <= 8'h2f;
		memory[16'h6eb] <= 8'hc9;
		memory[16'h6ec] <= 8'hdc;
		memory[16'h6ed] <= 8'hc4;
		memory[16'h6ee] <= 8'hc6;
		memory[16'h6ef] <= 8'h98;
		memory[16'h6f0] <= 8'h2c;
		memory[16'h6f1] <= 8'h11;
		memory[16'h6f2] <= 8'hf7;
		memory[16'h6f3] <= 8'h83;
		memory[16'h6f4] <= 8'hd6;
		memory[16'h6f5] <= 8'hee;
		memory[16'h6f6] <= 8'h3e;
		memory[16'h6f7] <= 8'hef;
		memory[16'h6f8] <= 8'h21;
		memory[16'h6f9] <= 8'h7e;
		memory[16'h6fa] <= 8'h95;
		memory[16'h6fb] <= 8'h99;
		memory[16'h6fc] <= 8'h36;
		memory[16'h6fd] <= 8'h53;
		memory[16'h6fe] <= 8'h85;
		memory[16'h6ff] <= 8'hee;
		memory[16'h700] <= 8'h7b;
		memory[16'h701] <= 8'hd6;
		memory[16'h702] <= 8'h2c;
		memory[16'h703] <= 8'hdb;
		memory[16'h704] <= 8'hfd;
		memory[16'h705] <= 8'h22;
		memory[16'h706] <= 8'h8c;
		memory[16'h707] <= 8'hc7;
		memory[16'h708] <= 8'hd3;
		memory[16'h709] <= 8'hbb;
		memory[16'h70a] <= 8'h90;
		memory[16'h70b] <= 8'hb0;
		memory[16'h70c] <= 8'h80;
		memory[16'h70d] <= 8'h56;
		memory[16'h70e] <= 8'h48;
		memory[16'h70f] <= 8'hac;
		memory[16'h710] <= 8'h68;
		memory[16'h711] <= 8'h3f;
		memory[16'h712] <= 8'h2f;
		memory[16'h713] <= 8'h3e;
		memory[16'h714] <= 8'h2d;
		memory[16'h715] <= 8'h6e;
		memory[16'h716] <= 8'h2d;
		memory[16'h717] <= 8'h4e;
		memory[16'h718] <= 8'hec;
		memory[16'h719] <= 8'hc2;
		memory[16'h71a] <= 8'he8;
		memory[16'h71b] <= 8'h22;
		memory[16'h71c] <= 8'h16;
		memory[16'h71d] <= 8'h6d;
		memory[16'h71e] <= 8'h11;
		memory[16'h71f] <= 8'h91;
		memory[16'h720] <= 8'h44;
		memory[16'h721] <= 8'h3d;
		memory[16'h722] <= 8'h6c;
		memory[16'h723] <= 8'h41;
		memory[16'h724] <= 8'h5f;
		memory[16'h725] <= 8'hf8;
		memory[16'h726] <= 8'h8;
		memory[16'h727] <= 8'h32;
		memory[16'h728] <= 8'hb4;
		memory[16'h729] <= 8'h99;
		memory[16'h72a] <= 8'he2;
		memory[16'h72b] <= 8'h34;
		memory[16'h72c] <= 8'hef;
		memory[16'h72d] <= 8'h2a;
		memory[16'h72e] <= 8'he0;
		memory[16'h72f] <= 8'h57;
		memory[16'h730] <= 8'h69;
		memory[16'h731] <= 8'h10;
		memory[16'h732] <= 8'h95;
		memory[16'h733] <= 8'h96;
		memory[16'h734] <= 8'h7e;
		memory[16'h735] <= 8'hc2;
		memory[16'h736] <= 8'he5;
		memory[16'h737] <= 8'h6a;
		memory[16'h738] <= 8'h85;
		memory[16'h739] <= 8'hcd;
		memory[16'h73a] <= 8'h8d;
		memory[16'h73b] <= 8'h9b;
		memory[16'h73c] <= 8'h3a;
		memory[16'h73d] <= 8'h9e;
		memory[16'h73e] <= 8'h2c;
		memory[16'h73f] <= 8'h7e;
		memory[16'h740] <= 8'hdb;
		memory[16'h741] <= 8'h99;
		memory[16'h742] <= 8'hc0;
		memory[16'h743] <= 8'h3a;
		memory[16'h744] <= 8'h91;
		memory[16'h745] <= 8'hc8;
		memory[16'h746] <= 8'h6c;
		memory[16'h747] <= 8'h45;
		memory[16'h748] <= 8'h61;
		memory[16'h749] <= 8'h4f;
		memory[16'h74a] <= 8'h79;
		memory[16'h74b] <= 8'h51;
		memory[16'h74c] <= 8'h79;
		memory[16'h74d] <= 8'h5a;
		memory[16'h74e] <= 8'ha8;
		memory[16'h74f] <= 8'he3;
		memory[16'h750] <= 8'h6a;
		memory[16'h751] <= 8'h3e;
		memory[16'h752] <= 8'h79;
		memory[16'h753] <= 8'he8;
		memory[16'h754] <= 8'h0;
		memory[16'h755] <= 8'h5e;
		memory[16'h756] <= 8'h52;
		memory[16'h757] <= 8'h85;
		memory[16'h758] <= 8'h2b;
		memory[16'h759] <= 8'hdf;
		memory[16'h75a] <= 8'h20;
		memory[16'h75b] <= 8'h66;
		memory[16'h75c] <= 8'h7d;
		memory[16'h75d] <= 8'h4d;
		memory[16'h75e] <= 8'he4;
		memory[16'h75f] <= 8'h58;
		memory[16'h760] <= 8'he6;
		memory[16'h761] <= 8'ha4;
		memory[16'h762] <= 8'h92;
		memory[16'h763] <= 8'h77;
		memory[16'h764] <= 8'h6d;
		memory[16'h765] <= 8'hff;
		memory[16'h766] <= 8'hbd;
		memory[16'h767] <= 8'hce;
		memory[16'h768] <= 8'h4e;
		memory[16'h769] <= 8'h36;
		memory[16'h76a] <= 8'h1f;
		memory[16'h76b] <= 8'hc7;
		memory[16'h76c] <= 8'h90;
		memory[16'h76d] <= 8'hc8;
		memory[16'h76e] <= 8'haa;
		memory[16'h76f] <= 8'hfa;
		memory[16'h770] <= 8'h6;
		memory[16'h771] <= 8'h24;
		memory[16'h772] <= 8'he2;
		memory[16'h773] <= 8'h6;
		memory[16'h774] <= 8'h82;
		memory[16'h775] <= 8'h35;
		memory[16'h776] <= 8'h8c;
		memory[16'h777] <= 8'hae;
		memory[16'h778] <= 8'h14;
		memory[16'h779] <= 8'hac;
		memory[16'h77a] <= 8'h14;
		memory[16'h77b] <= 8'h92;
		memory[16'h77c] <= 8'hf9;
		memory[16'h77d] <= 8'hf8;
		memory[16'h77e] <= 8'hea;
		memory[16'h77f] <= 8'hdf;
		memory[16'h780] <= 8'h9d;
		memory[16'h781] <= 8'h7d;
		memory[16'h782] <= 8'h57;
		memory[16'h783] <= 8'ha;
		memory[16'h784] <= 8'h7c;
		memory[16'h785] <= 8'h14;
		memory[16'h786] <= 8'hd8;
		memory[16'h787] <= 8'hca;
		memory[16'h788] <= 8'h4a;
		memory[16'h789] <= 8'hf8;
		memory[16'h78a] <= 8'h91;
		memory[16'h78b] <= 8'hdb;
		memory[16'h78c] <= 8'hc0;
		memory[16'h78d] <= 8'h3c;
		memory[16'h78e] <= 8'hd5;
		memory[16'h78f] <= 8'hc6;
		memory[16'h790] <= 8'h60;
		memory[16'h791] <= 8'hb8;
		memory[16'h792] <= 8'hcc;
		memory[16'h793] <= 8'he2;
		memory[16'h794] <= 8'hed;
		memory[16'h795] <= 8'h58;
		memory[16'h796] <= 8'h90;
		memory[16'h797] <= 8'h1;
		memory[16'h798] <= 8'h5;
		memory[16'h799] <= 8'ha4;
		memory[16'h79a] <= 8'h93;
		memory[16'h79b] <= 8'hfe;
		memory[16'h79c] <= 8'h9d;
		memory[16'h79d] <= 8'h7e;
		memory[16'h79e] <= 8'hde;
		memory[16'h79f] <= 8'h3a;
		memory[16'h7a0] <= 8'hfb;
		memory[16'h7a1] <= 8'h35;
		memory[16'h7a2] <= 8'h44;
		memory[16'h7a3] <= 8'h77;
		memory[16'h7a4] <= 8'h49;
		memory[16'h7a5] <= 8'h1c;
		memory[16'h7a6] <= 8'h41;
		memory[16'h7a7] <= 8'h93;
		memory[16'h7a8] <= 8'h14;
		memory[16'h7a9] <= 8'hd2;
		memory[16'h7aa] <= 8'h6e;
		memory[16'h7ab] <= 8'hd4;
		memory[16'h7ac] <= 8'he;
		memory[16'h7ad] <= 8'h44;
		memory[16'h7ae] <= 8'h9a;
		memory[16'h7af] <= 8'h6e;
		memory[16'h7b0] <= 8'hfc;
		memory[16'h7b1] <= 8'h67;
		memory[16'h7b2] <= 8'h51;
		memory[16'h7b3] <= 8'he9;
		memory[16'h7b4] <= 8'hbf;
		memory[16'h7b5] <= 8'he1;
		memory[16'h7b6] <= 8'hea;
		memory[16'h7b7] <= 8'hc4;
		memory[16'h7b8] <= 8'h86;
		memory[16'h7b9] <= 8'h7e;
		memory[16'h7ba] <= 8'hc3;
		memory[16'h7bb] <= 8'h23;
		memory[16'h7bc] <= 8'hfc;
		memory[16'h7bd] <= 8'ha1;
		memory[16'h7be] <= 8'h5d;
		memory[16'h7bf] <= 8'hf7;
		memory[16'h7c0] <= 8'hd6;
		memory[16'h7c1] <= 8'ha1;
		memory[16'h7c2] <= 8'h6e;
		memory[16'h7c3] <= 8'h1f;
		memory[16'h7c4] <= 8'hbd;
		memory[16'h7c5] <= 8'haf;
		memory[16'h7c6] <= 8'hb2;
		memory[16'h7c7] <= 8'hd2;
		memory[16'h7c8] <= 8'h81;
		memory[16'h7c9] <= 8'h21;
		memory[16'h7ca] <= 8'ha6;
		memory[16'h7cb] <= 8'h90;
		memory[16'h7cc] <= 8'h65;
		memory[16'h7cd] <= 8'h41;
		memory[16'h7ce] <= 8'hfe;
		memory[16'h7cf] <= 8'h61;
		memory[16'h7d0] <= 8'ha8;
		memory[16'h7d1] <= 8'h4f;
		memory[16'h7d2] <= 8'h4a;
		memory[16'h7d3] <= 8'h67;
		memory[16'h7d4] <= 8'h31;
		memory[16'h7d5] <= 8'h34;
		memory[16'h7d6] <= 8'h2c;
		memory[16'h7d7] <= 8'hb7;
		memory[16'h7d8] <= 8'hb2;
		memory[16'h7d9] <= 8'hef;
		memory[16'h7da] <= 8'hda;
		memory[16'h7db] <= 8'hae;
		memory[16'h7dc] <= 8'h90;
		memory[16'h7dd] <= 8'h37;
		memory[16'h7de] <= 8'ha5;
		memory[16'h7df] <= 8'h66;
		memory[16'h7e0] <= 8'hd8;
		memory[16'h7e1] <= 8'h13;
		memory[16'h7e2] <= 8'h85;
		memory[16'h7e3] <= 8'h95;
		memory[16'h7e4] <= 8'hc2;
		memory[16'h7e5] <= 8'h37;
		memory[16'h7e6] <= 8'h67;
		memory[16'h7e7] <= 8'h44;
		memory[16'h7e8] <= 8'h58;
		memory[16'h7e9] <= 8'he;
		memory[16'h7ea] <= 8'hd4;
		memory[16'h7eb] <= 8'hbd;
		memory[16'h7ec] <= 8'h4f;
		memory[16'h7ed] <= 8'hd2;
		memory[16'h7ee] <= 8'h1e;
		memory[16'h7ef] <= 8'hf7;
		memory[16'h7f0] <= 8'h22;
		memory[16'h7f1] <= 8'h68;
		memory[16'h7f2] <= 8'h5e;
		memory[16'h7f3] <= 8'h53;
		memory[16'h7f4] <= 8'h9d;
		memory[16'h7f5] <= 8'h8a;
		memory[16'h7f6] <= 8'ha;
		memory[16'h7f7] <= 8'h4f;
		memory[16'h7f8] <= 8'h79;
		memory[16'h7f9] <= 8'he4;
		memory[16'h7fa] <= 8'hfe;
		memory[16'h7fb] <= 8'h9;
		memory[16'h7fc] <= 8'h1b;
		memory[16'h7fd] <= 8'ha3;
		memory[16'h7fe] <= 8'h6f;
		memory[16'h7ff] <= 8'hf3;
		memory[16'h800] <= 8'hb7;
		memory[16'h801] <= 8'hf4;
		memory[16'h802] <= 8'h88;
		memory[16'h803] <= 8'h79;
		memory[16'h804] <= 8'h2c;
		memory[16'h805] <= 8'hf0;
		memory[16'h806] <= 8'hbd;
		memory[16'h807] <= 8'h84;
		memory[16'h808] <= 8'hfe;
		memory[16'h809] <= 8'h91;
		memory[16'h80a] <= 8'h42;
		memory[16'h80b] <= 8'h4d;
		memory[16'h80c] <= 8'h64;
		memory[16'h80d] <= 8'h60;
		memory[16'h80e] <= 8'h44;
		memory[16'h80f] <= 8'h86;
		memory[16'h810] <= 8'hc9;
		memory[16'h811] <= 8'ha2;
		memory[16'h812] <= 8'hd9;
		memory[16'h813] <= 8'h66;
		memory[16'h814] <= 8'h2d;
		memory[16'h815] <= 8'he3;
		memory[16'h816] <= 8'hb5;
		memory[16'h817] <= 8'ha6;
		memory[16'h818] <= 8'hc7;
		memory[16'h819] <= 8'hb3;
		memory[16'h81a] <= 8'hb0;
		memory[16'h81b] <= 8'he2;
		memory[16'h81c] <= 8'h57;
		memory[16'h81d] <= 8'h1f;
		memory[16'h81e] <= 8'hd5;
		memory[16'h81f] <= 8'he;
		memory[16'h820] <= 8'h14;
		memory[16'h821] <= 8'h5d;
		memory[16'h822] <= 8'h87;
		memory[16'h823] <= 8'h40;
		memory[16'h824] <= 8'h4d;
		memory[16'h825] <= 8'h45;
		memory[16'h826] <= 8'hc4;
		memory[16'h827] <= 8'h4b;
		memory[16'h828] <= 8'hd6;
		memory[16'h829] <= 8'h6;
		memory[16'h82a] <= 8'h98;
		memory[16'h82b] <= 8'h3a;
		memory[16'h82c] <= 8'h67;
		memory[16'h82d] <= 8'hdc;
		memory[16'h82e] <= 8'hc0;
		memory[16'h82f] <= 8'h30;
		memory[16'h830] <= 8'h7f;
		memory[16'h831] <= 8'h99;
		memory[16'h832] <= 8'h96;
		memory[16'h833] <= 8'hac;
		memory[16'h834] <= 8'h7c;
		memory[16'h835] <= 8'h4b;
		memory[16'h836] <= 8'h52;
		memory[16'h837] <= 8'h43;
		memory[16'h838] <= 8'hff;
		memory[16'h839] <= 8'h2;
		memory[16'h83a] <= 8'h25;
		memory[16'h83b] <= 8'h56;
		memory[16'h83c] <= 8'h22;
		memory[16'h83d] <= 8'hfa;
		memory[16'h83e] <= 8'h64;
		memory[16'h83f] <= 8'h36;
		memory[16'h840] <= 8'h58;
		memory[16'h841] <= 8'heb;
		memory[16'h842] <= 8'h76;
		memory[16'h843] <= 8'ha5;
		memory[16'h844] <= 8'h30;
		memory[16'h845] <= 8'h3a;
		memory[16'h846] <= 8'hf1;
		memory[16'h847] <= 8'h7;
		memory[16'h848] <= 8'h41;
		memory[16'h849] <= 8'h89;
		memory[16'h84a] <= 8'h41;
		memory[16'h84b] <= 8'ha8;
		memory[16'h84c] <= 8'h66;
		memory[16'h84d] <= 8'h2;
		memory[16'h84e] <= 8'hd8;
		memory[16'h84f] <= 8'he5;
		memory[16'h850] <= 8'h9b;
		memory[16'h851] <= 8'h6e;
		memory[16'h852] <= 8'h91;
		memory[16'h853] <= 8'h18;
		memory[16'h854] <= 8'hb9;
		memory[16'h855] <= 8'he3;
		memory[16'h856] <= 8'h5b;
		memory[16'h857] <= 8'hb8;
		memory[16'h858] <= 8'he6;
		memory[16'h859] <= 8'h81;
		memory[16'h85a] <= 8'he;
		memory[16'h85b] <= 8'h8;
		memory[16'h85c] <= 8'h7b;
		memory[16'h85d] <= 8'h72;
		memory[16'h85e] <= 8'h3e;
		memory[16'h85f] <= 8'hd3;
		memory[16'h860] <= 8'h5e;
		memory[16'h861] <= 8'hb4;
		memory[16'h862] <= 8'h79;
		memory[16'h863] <= 8'h8e;
		memory[16'h864] <= 8'hee;
		memory[16'h865] <= 8'h6a;
		memory[16'h866] <= 8'h95;
		memory[16'h867] <= 8'h2f;
		memory[16'h868] <= 8'hf3;
		memory[16'h869] <= 8'hd7;
		memory[16'h86a] <= 8'hd7;
		memory[16'h86b] <= 8'h59;
		memory[16'h86c] <= 8'hd9;
		memory[16'h86d] <= 8'haf;
		memory[16'h86e] <= 8'h3e;
		memory[16'h86f] <= 8'h74;
		memory[16'h870] <= 8'h1d;
		memory[16'h871] <= 8'hcf;
		memory[16'h872] <= 8'h8c;
		memory[16'h873] <= 8'hd7;
		memory[16'h874] <= 8'hb3;
		memory[16'h875] <= 8'he8;
		memory[16'h876] <= 8'h8f;
		memory[16'h877] <= 8'h99;
		memory[16'h878] <= 8'h69;
		memory[16'h879] <= 8'h9e;
		memory[16'h87a] <= 8'ha1;
		memory[16'h87b] <= 8'he4;
		memory[16'h87c] <= 8'h10;
		memory[16'h87d] <= 8'hdf;
		memory[16'h87e] <= 8'hb8;
		memory[16'h87f] <= 8'h6e;
		memory[16'h880] <= 8'h93;
		memory[16'h881] <= 8'h31;
		memory[16'h882] <= 8'hfd;
		memory[16'h883] <= 8'h81;
		memory[16'h884] <= 8'h9b;
		memory[16'h885] <= 8'h92;
		memory[16'h886] <= 8'hb1;
		memory[16'h887] <= 8'h8e;
		memory[16'h888] <= 8'h69;
		memory[16'h889] <= 8'h88;
		memory[16'h88a] <= 8'he8;
		memory[16'h88b] <= 8'h42;
		memory[16'h88c] <= 8'h38;
		memory[16'h88d] <= 8'h26;
		memory[16'h88e] <= 8'hb7;
		memory[16'h88f] <= 8'h55;
		memory[16'h890] <= 8'hf6;
		memory[16'h891] <= 8'h43;
		memory[16'h892] <= 8'h2c;
		memory[16'h893] <= 8'ha9;
		memory[16'h894] <= 8'h2b;
		memory[16'h895] <= 8'hbc;
		memory[16'h896] <= 8'h42;
		memory[16'h897] <= 8'h94;
		memory[16'h898] <= 8'h5a;
		memory[16'h899] <= 8'he3;
		memory[16'h89a] <= 8'h79;
		memory[16'h89b] <= 8'h6a;
		memory[16'h89c] <= 8'hc2;
		memory[16'h89d] <= 8'h31;
		memory[16'h89e] <= 8'hd9;
		memory[16'h89f] <= 8'h55;
		memory[16'h8a0] <= 8'h62;
		memory[16'h8a1] <= 8'hd6;
		memory[16'h8a2] <= 8'hd6;
		memory[16'h8a3] <= 8'hfd;
		memory[16'h8a4] <= 8'h68;
		memory[16'h8a5] <= 8'h87;
		memory[16'h8a6] <= 8'h8b;
		memory[16'h8a7] <= 8'hd2;
		memory[16'h8a8] <= 8'h10;
		memory[16'h8a9] <= 8'h73;
		memory[16'h8aa] <= 8'h14;
		memory[16'h8ab] <= 8'h48;
		memory[16'h8ac] <= 8'h9a;
		memory[16'h8ad] <= 8'hcb;
		memory[16'h8ae] <= 8'h9d;
		memory[16'h8af] <= 8'h90;
		memory[16'h8b0] <= 8'hf;
		memory[16'h8b1] <= 8'hca;
		memory[16'h8b2] <= 8'h39;
		memory[16'h8b3] <= 8'h3a;
		memory[16'h8b4] <= 8'h86;
		memory[16'h8b5] <= 8'h7b;
		memory[16'h8b6] <= 8'hcf;
		memory[16'h8b7] <= 8'he0;
		memory[16'h8b8] <= 8'h5e;
		memory[16'h8b9] <= 8'h48;
		memory[16'h8ba] <= 8'h4a;
		memory[16'h8bb] <= 8'h20;
		memory[16'h8bc] <= 8'h79;
		memory[16'h8bd] <= 8'h23;
		memory[16'h8be] <= 8'h75;
		memory[16'h8bf] <= 8'hdb;
		memory[16'h8c0] <= 8'hf9;
		memory[16'h8c1] <= 8'h4b;
		memory[16'h8c2] <= 8'hd8;
		memory[16'h8c3] <= 8'h62;
		memory[16'h8c4] <= 8'hd3;
		memory[16'h8c5] <= 8'h63;
		memory[16'h8c6] <= 8'h34;
		memory[16'h8c7] <= 8'he3;
		memory[16'h8c8] <= 8'hd7;
		memory[16'h8c9] <= 8'h48;
		memory[16'h8ca] <= 8'h2b;
		memory[16'h8cb] <= 8'h71;
		memory[16'h8cc] <= 8'h14;
		memory[16'h8cd] <= 8'hc8;
		memory[16'h8ce] <= 8'h1;
		memory[16'h8cf] <= 8'h23;
		memory[16'h8d0] <= 8'h92;
		memory[16'h8d1] <= 8'h3a;
		memory[16'h8d2] <= 8'h5d;
		memory[16'h8d3] <= 8'h18;
		memory[16'h8d4] <= 8'hb5;
		memory[16'h8d5] <= 8'h2c;
		memory[16'h8d6] <= 8'hf8;
		memory[16'h8d7] <= 8'h13;
		memory[16'h8d8] <= 8'h74;
		memory[16'h8d9] <= 8'h43;
		memory[16'h8da] <= 8'h33;
		memory[16'h8db] <= 8'hed;
		memory[16'h8dc] <= 8'h66;
		memory[16'h8dd] <= 8'ha8;
		memory[16'h8de] <= 8'hc8;
		memory[16'h8df] <= 8'h60;
		memory[16'h8e0] <= 8'hf3;
		memory[16'h8e1] <= 8'ha0;
		memory[16'h8e2] <= 8'hc2;
		memory[16'h8e3] <= 8'hc6;
		memory[16'h8e4] <= 8'h4;
		memory[16'h8e5] <= 8'hf6;
		memory[16'h8e6] <= 8'ha9;
		memory[16'h8e7] <= 8'hdb;
		memory[16'h8e8] <= 8'h3e;
		memory[16'h8e9] <= 8'hd4;
		memory[16'h8ea] <= 8'h4c;
		memory[16'h8eb] <= 8'h52;
		memory[16'h8ec] <= 8'h9d;
		memory[16'h8ed] <= 8'h4d;
		memory[16'h8ee] <= 8'h75;
		memory[16'h8ef] <= 8'h2f;
		memory[16'h8f0] <= 8'h87;
		memory[16'h8f1] <= 8'hd3;
		memory[16'h8f2] <= 8'h48;
		memory[16'h8f3] <= 8'h3c;
		memory[16'h8f4] <= 8'hff;
		memory[16'h8f5] <= 8'h40;
		memory[16'h8f6] <= 8'h4f;
		memory[16'h8f7] <= 8'h74;
		memory[16'h8f8] <= 8'h83;
		memory[16'h8f9] <= 8'h82;
		memory[16'h8fa] <= 8'h61;
		memory[16'h8fb] <= 8'hea;
		memory[16'h8fc] <= 8'h2a;
		memory[16'h8fd] <= 8'h2a;
		memory[16'h8fe] <= 8'h4a;
		memory[16'h8ff] <= 8'h1d;
		memory[16'h900] <= 8'hca;
		memory[16'h901] <= 8'hc;
		memory[16'h902] <= 8'he4;
		memory[16'h903] <= 8'hce;
		memory[16'h904] <= 8'h2;
		memory[16'h905] <= 8'h8d;
		memory[16'h906] <= 8'ha9;
		memory[16'h907] <= 8'h40;
		memory[16'h908] <= 8'h62;
		memory[16'h909] <= 8'hf5;
		memory[16'h90a] <= 8'h93;
		memory[16'h90b] <= 8'hff;
		memory[16'h90c] <= 8'h42;
		memory[16'h90d] <= 8'h8;
		memory[16'h90e] <= 8'h2e;
		memory[16'h90f] <= 8'hc9;
		memory[16'h910] <= 8'hdb;
		memory[16'h911] <= 8'h76;
		memory[16'h912] <= 8'h5;
		memory[16'h913] <= 8'hdb;
		memory[16'h914] <= 8'hb7;
		memory[16'h915] <= 8'h54;
		memory[16'h916] <= 8'h4f;
		memory[16'h917] <= 8'h3a;
		memory[16'h918] <= 8'hd6;
		memory[16'h919] <= 8'hb0;
		memory[16'h91a] <= 8'h24;
		memory[16'h91b] <= 8'h0;
		memory[16'h91c] <= 8'hda;
		memory[16'h91d] <= 8'h6e;
		memory[16'h91e] <= 8'h1e;
		memory[16'h91f] <= 8'ha5;
		memory[16'h920] <= 8'h7a;
		memory[16'h921] <= 8'h2;
		memory[16'h922] <= 8'h73;
		memory[16'h923] <= 8'h7c;
		memory[16'h924] <= 8'h8f;
		memory[16'h925] <= 8'h1d;
		memory[16'h926] <= 8'hbd;
		memory[16'h927] <= 8'hf1;
		memory[16'h928] <= 8'h12;
		memory[16'h929] <= 8'h50;
		memory[16'h92a] <= 8'hf0;
		memory[16'h92b] <= 8'h55;
		memory[16'h92c] <= 8'h58;
		memory[16'h92d] <= 8'h1f;
		memory[16'h92e] <= 8'h1e;
		memory[16'h92f] <= 8'h34;
		memory[16'h930] <= 8'h95;
		memory[16'h931] <= 8'h24;
		memory[16'h932] <= 8'hf;
		memory[16'h933] <= 8'h4c;
		memory[16'h934] <= 8'h78;
		memory[16'h935] <= 8'h5e;
		memory[16'h936] <= 8'h87;
		memory[16'h937] <= 8'h4f;
		memory[16'h938] <= 8'he;
		memory[16'h939] <= 8'hab;
		memory[16'h93a] <= 8'h4f;
		memory[16'h93b] <= 8'he9;
		memory[16'h93c] <= 8'h1a;
		memory[16'h93d] <= 8'h6d;
		memory[16'h93e] <= 8'h8e;
		memory[16'h93f] <= 8'h94;
		memory[16'h940] <= 8'h6f;
		memory[16'h941] <= 8'h1;
		memory[16'h942] <= 8'h11;
		memory[16'h943] <= 8'hff;
		memory[16'h944] <= 8'h1e;
		memory[16'h945] <= 8'hce;
		memory[16'h946] <= 8'hf0;
		memory[16'h947] <= 8'h31;
		memory[16'h948] <= 8'h1e;
		memory[16'h949] <= 8'he1;
		memory[16'h94a] <= 8'h86;
		memory[16'h94b] <= 8'h76;
		memory[16'h94c] <= 8'h0;
		memory[16'h94d] <= 8'ha4;
		memory[16'h94e] <= 8'haa;
		memory[16'h94f] <= 8'h95;
		memory[16'h950] <= 8'hc8;
		memory[16'h951] <= 8'hb9;
		memory[16'h952] <= 8'he2;
		memory[16'h953] <= 8'h41;
		memory[16'h954] <= 8'h17;
		memory[16'h955] <= 8'h69;
		memory[16'h956] <= 8'h90;
		memory[16'h957] <= 8'h26;
		memory[16'h958] <= 8'h14;
		memory[16'h959] <= 8'hdf;
		memory[16'h95a] <= 8'hf;
		memory[16'h95b] <= 8'h2e;
		memory[16'h95c] <= 8'h4d;
		memory[16'h95d] <= 8'h9d;
		memory[16'h95e] <= 8'hc3;
		memory[16'h95f] <= 8'hbc;
		memory[16'h960] <= 8'h9e;
		memory[16'h961] <= 8'hd4;
		memory[16'h962] <= 8'hbb;
		memory[16'h963] <= 8'hbd;
		memory[16'h964] <= 8'ha2;
		memory[16'h965] <= 8'hac;
		memory[16'h966] <= 8'hee;
		memory[16'h967] <= 8'hc0;
		memory[16'h968] <= 8'h8d;
		memory[16'h969] <= 8'h74;
		memory[16'h96a] <= 8'h36;
		memory[16'h96b] <= 8'h8d;
		memory[16'h96c] <= 8'h18;
		memory[16'h96d] <= 8'he1;
		memory[16'h96e] <= 8'h22;
		memory[16'h96f] <= 8'he1;
		memory[16'h970] <= 8'h9a;
		memory[16'h971] <= 8'h4;
		memory[16'h972] <= 8'h22;
		memory[16'h973] <= 8'hb2;
		memory[16'h974] <= 8'h6d;
		memory[16'h975] <= 8'hb2;
		memory[16'h976] <= 8'hd8;
		memory[16'h977] <= 8'h82;
		memory[16'h978] <= 8'h91;
		memory[16'h979] <= 8'he7;
		memory[16'h97a] <= 8'hb0;
		memory[16'h97b] <= 8'hde;
		memory[16'h97c] <= 8'h84;
		memory[16'h97d] <= 8'h73;
		memory[16'h97e] <= 8'h9b;
		memory[16'h97f] <= 8'h22;
		memory[16'h980] <= 8'h47;
		memory[16'h981] <= 8'h56;
		memory[16'h982] <= 8'hdf;
		memory[16'h983] <= 8'he9;
		memory[16'h984] <= 8'h2;
		memory[16'h985] <= 8'hcd;
		memory[16'h986] <= 8'ha9;
		memory[16'h987] <= 8'h8f;
		memory[16'h988] <= 8'h41;
		memory[16'h989] <= 8'he0;
		memory[16'h98a] <= 8'h1c;
		memory[16'h98b] <= 8'h5a;
		memory[16'h98c] <= 8'hc1;
		memory[16'h98d] <= 8'h3f;
		memory[16'h98e] <= 8'h3b;
		memory[16'h98f] <= 8'h5b;
		memory[16'h990] <= 8'h43;
		memory[16'h991] <= 8'h5d;
		memory[16'h992] <= 8'hd;
		memory[16'h993] <= 8'hb1;
		memory[16'h994] <= 8'hf;
		memory[16'h995] <= 8'he5;
		memory[16'h996] <= 8'h33;
		memory[16'h997] <= 8'ha0;
		memory[16'h998] <= 8'hcc;
		memory[16'h999] <= 8'he3;
		memory[16'h99a] <= 8'h7f;
		memory[16'h99b] <= 8'h50;
		memory[16'h99c] <= 8'h57;
		memory[16'h99d] <= 8'h1a;
		memory[16'h99e] <= 8'h73;
		memory[16'h99f] <= 8'h9e;
		memory[16'h9a0] <= 8'h70;
		memory[16'h9a1] <= 8'h52;
		memory[16'h9a2] <= 8'h88;
		memory[16'h9a3] <= 8'h73;
		memory[16'h9a4] <= 8'h20;
		memory[16'h9a5] <= 8'h31;
		memory[16'h9a6] <= 8'h2;
		memory[16'h9a7] <= 8'h61;
		memory[16'h9a8] <= 8'h11;
		memory[16'h9a9] <= 8'h1f;
		memory[16'h9aa] <= 8'hbb;
		memory[16'h9ab] <= 8'hd2;
		memory[16'h9ac] <= 8'h5e;
		memory[16'h9ad] <= 8'hf6;
		memory[16'h9ae] <= 8'h2e;
		memory[16'h9af] <= 8'ha1;
		memory[16'h9b0] <= 8'h53;
		memory[16'h9b1] <= 8'h3b;
		memory[16'h9b2] <= 8'h52;
		memory[16'h9b3] <= 8'h62;
		memory[16'h9b4] <= 8'h21;
		memory[16'h9b5] <= 8'h85;
		memory[16'h9b6] <= 8'h3;
		memory[16'h9b7] <= 8'hed;
		memory[16'h9b8] <= 8'h69;
		memory[16'h9b9] <= 8'h82;
		memory[16'h9ba] <= 8'h3e;
		memory[16'h9bb] <= 8'hc0;
		memory[16'h9bc] <= 8'h9c;
		memory[16'h9bd] <= 8'hb1;
		memory[16'h9be] <= 8'h5e;
		memory[16'h9bf] <= 8'hc;
		memory[16'h9c0] <= 8'h3;
		memory[16'h9c1] <= 8'he6;
		memory[16'h9c2] <= 8'h7f;
		memory[16'h9c3] <= 8'h23;
		memory[16'h9c4] <= 8'h18;
		memory[16'h9c5] <= 8'h82;
		memory[16'h9c6] <= 8'h85;
		memory[16'h9c7] <= 8'h29;
		memory[16'h9c8] <= 8'ha1;
		memory[16'h9c9] <= 8'h40;
		memory[16'h9ca] <= 8'hfc;
		memory[16'h9cb] <= 8'hff;
		memory[16'h9cc] <= 8'h37;
		memory[16'h9cd] <= 8'h2a;
		memory[16'h9ce] <= 8'ha0;
		memory[16'h9cf] <= 8'h8a;
		memory[16'h9d0] <= 8'h65;
		memory[16'h9d1] <= 8'hf3;
		memory[16'h9d2] <= 8'hed;
		memory[16'h9d3] <= 8'h86;
		memory[16'h9d4] <= 8'h78;
		memory[16'h9d5] <= 8'hf0;
		memory[16'h9d6] <= 8'h74;
		memory[16'h9d7] <= 8'he1;
		memory[16'h9d8] <= 8'h72;
		memory[16'h9d9] <= 8'hb2;
		memory[16'h9da] <= 8'ha1;
		memory[16'h9db] <= 8'he;
		memory[16'h9dc] <= 8'h63;
		memory[16'h9dd] <= 8'h0;
		memory[16'h9de] <= 8'h1a;
		memory[16'h9df] <= 8'h66;
		memory[16'h9e0] <= 8'he6;
		memory[16'h9e1] <= 8'h9a;
		memory[16'h9e2] <= 8'h8a;
		memory[16'h9e3] <= 8'hfe;
		memory[16'h9e4] <= 8'h1c;
		memory[16'h9e5] <= 8'hf;
		memory[16'h9e6] <= 8'h28;
		memory[16'h9e7] <= 8'hbd;
		memory[16'h9e8] <= 8'h4f;
		memory[16'h9e9] <= 8'h24;
		memory[16'h9ea] <= 8'hbc;
		memory[16'h9eb] <= 8'h86;
		memory[16'h9ec] <= 8'h4e;
		memory[16'h9ed] <= 8'h5c;
		memory[16'h9ee] <= 8'h11;
		memory[16'h9ef] <= 8'hb3;
		memory[16'h9f0] <= 8'h4f;
		memory[16'h9f1] <= 8'hfe;
		memory[16'h9f2] <= 8'h3a;
		memory[16'h9f3] <= 8'hc8;
		memory[16'h9f4] <= 8'hee;
		memory[16'h9f5] <= 8'hae;
		memory[16'h9f6] <= 8'ha9;
		memory[16'h9f7] <= 8'h60;
		memory[16'h9f8] <= 8'h60;
		memory[16'h9f9] <= 8'h4b;
		memory[16'h9fa] <= 8'h6e;
		memory[16'h9fb] <= 8'hc3;
		memory[16'h9fc] <= 8'h4b;
		memory[16'h9fd] <= 8'h88;
		memory[16'h9fe] <= 8'h29;
		memory[16'h9ff] <= 8'h31;
		memory[16'ha00] <= 8'h22;
		memory[16'ha01] <= 8'hb3;
		memory[16'ha02] <= 8'h30;
		memory[16'ha03] <= 8'h3e;
		memory[16'ha04] <= 8'hc2;
		memory[16'ha05] <= 8'h58;
		memory[16'ha06] <= 8'hfb;
		memory[16'ha07] <= 8'h12;
		memory[16'ha08] <= 8'h7c;
		memory[16'ha09] <= 8'hb7;
		memory[16'ha0a] <= 8'h98;
		memory[16'ha0b] <= 8'hca;
		memory[16'ha0c] <= 8'h14;
		memory[16'ha0d] <= 8'ha9;
		memory[16'ha0e] <= 8'h7d;
		memory[16'ha0f] <= 8'h63;
		memory[16'ha10] <= 8'ha7;
		memory[16'ha11] <= 8'hb7;
		memory[16'ha12] <= 8'h2b;
		memory[16'ha13] <= 8'h95;
		memory[16'ha14] <= 8'h65;
		memory[16'ha15] <= 8'hd5;
		memory[16'ha16] <= 8'hf5;
		memory[16'ha17] <= 8'hc5;
		memory[16'ha18] <= 8'h20;
		memory[16'ha19] <= 8'h63;
		memory[16'ha1a] <= 8'h88;
		memory[16'ha1b] <= 8'h6b;
		memory[16'ha1c] <= 8'hec;
		memory[16'ha1d] <= 8'hb2;
		memory[16'ha1e] <= 8'h9c;
		memory[16'ha1f] <= 8'he;
		memory[16'ha20] <= 8'h65;
		memory[16'ha21] <= 8'hcc;
		memory[16'ha22] <= 8'h4d;
		memory[16'ha23] <= 8'h28;
		memory[16'ha24] <= 8'h24;
		memory[16'ha25] <= 8'h48;
		memory[16'ha26] <= 8'h3a;
		memory[16'ha27] <= 8'ha0;
		memory[16'ha28] <= 8'h0;
		memory[16'ha29] <= 8'hd2;
		memory[16'ha2a] <= 8'h6a;
		memory[16'ha2b] <= 8'h14;
		memory[16'ha2c] <= 8'h7c;
		memory[16'ha2d] <= 8'he8;
		memory[16'ha2e] <= 8'h77;
		memory[16'ha2f] <= 8'h23;
		memory[16'ha30] <= 8'h9f;
		memory[16'ha31] <= 8'ha3;
		memory[16'ha32] <= 8'hb9;
		memory[16'ha33] <= 8'h5;
		memory[16'ha34] <= 8'h78;
		memory[16'ha35] <= 8'hae;
		memory[16'ha36] <= 8'hca;
		memory[16'ha37] <= 8'h98;
		memory[16'ha38] <= 8'h12;
		memory[16'ha39] <= 8'h53;
		memory[16'ha3a] <= 8'h3;
		memory[16'ha3b] <= 8'hfe;
		memory[16'ha3c] <= 8'h5;
		memory[16'ha3d] <= 8'h9f;
		memory[16'ha3e] <= 8'hc;
		memory[16'ha3f] <= 8'h6a;
		memory[16'ha40] <= 8'h6c;
		memory[16'ha41] <= 8'h59;
		memory[16'ha42] <= 8'h92;
		memory[16'ha43] <= 8'h90;
		memory[16'ha44] <= 8'ha2;
		memory[16'ha45] <= 8'hcc;
		memory[16'ha46] <= 8'h31;
		memory[16'ha47] <= 8'ha2;
		memory[16'ha48] <= 8'h9f;
		memory[16'ha49] <= 8'h9b;
		memory[16'ha4a] <= 8'hb6;
		memory[16'ha4b] <= 8'h1b;
		memory[16'ha4c] <= 8'h83;
		memory[16'ha4d] <= 8'h2d;
		memory[16'ha4e] <= 8'h3e;
		memory[16'ha4f] <= 8'h23;
		memory[16'ha50] <= 8'hd0;
		memory[16'ha51] <= 8'hf7;
		memory[16'ha52] <= 8'h28;
		memory[16'ha53] <= 8'h48;
		memory[16'ha54] <= 8'ha6;
		memory[16'ha55] <= 8'hf2;
		memory[16'ha56] <= 8'he0;
		memory[16'ha57] <= 8'hb8;
		memory[16'ha58] <= 8'h45;
		memory[16'ha59] <= 8'he3;
		memory[16'ha5a] <= 8'hb6;
		memory[16'ha5b] <= 8'h4a;
		memory[16'ha5c] <= 8'h83;
		memory[16'ha5d] <= 8'hc2;
		memory[16'ha5e] <= 8'hb5;
		memory[16'ha5f] <= 8'hef;
		memory[16'ha60] <= 8'h1c;
		memory[16'ha61] <= 8'h47;
		memory[16'ha62] <= 8'h7f;
		memory[16'ha63] <= 8'hbe;
		memory[16'ha64] <= 8'h14;
		memory[16'ha65] <= 8'hb0;
		memory[16'ha66] <= 8'h60;
		memory[16'ha67] <= 8'hb3;
		memory[16'ha68] <= 8'h4c;
		memory[16'ha69] <= 8'h16;
		memory[16'ha6a] <= 8'hce;
		memory[16'ha6b] <= 8'hcf;
		memory[16'ha6c] <= 8'h43;
		memory[16'ha6d] <= 8'hc;
		memory[16'ha6e] <= 8'hf2;
		memory[16'ha6f] <= 8'h14;
		memory[16'ha70] <= 8'h4;
		memory[16'ha71] <= 8'h1a;
		memory[16'ha72] <= 8'h5c;
		memory[16'ha73] <= 8'haa;
		memory[16'ha74] <= 8'hd;
		memory[16'ha75] <= 8'h3d;
		memory[16'ha76] <= 8'h62;
		memory[16'ha77] <= 8'h52;
		memory[16'ha78] <= 8'h20;
		memory[16'ha79] <= 8'h18;
		memory[16'ha7a] <= 8'h9d;
		memory[16'ha7b] <= 8'ha3;
		memory[16'ha7c] <= 8'hda;
		memory[16'ha7d] <= 8'h52;
		memory[16'ha7e] <= 8'h92;
		memory[16'ha7f] <= 8'hf6;
		memory[16'ha80] <= 8'h99;
		memory[16'ha81] <= 8'h12;
		memory[16'ha82] <= 8'hb4;
		memory[16'ha83] <= 8'had;
		memory[16'ha84] <= 8'hc2;
		memory[16'ha85] <= 8'h14;
		memory[16'ha86] <= 8'h60;
		memory[16'ha87] <= 8'he;
		memory[16'ha88] <= 8'h2a;
		memory[16'ha89] <= 8'h2e;
		memory[16'ha8a] <= 8'hde;
		memory[16'ha8b] <= 8'h6e;
		memory[16'ha8c] <= 8'h3b;
		memory[16'ha8d] <= 8'hd0;
		memory[16'ha8e] <= 8'h82;
		memory[16'ha8f] <= 8'h3f;
		memory[16'ha90] <= 8'heb;
		memory[16'ha91] <= 8'hde;
		memory[16'ha92] <= 8'he9;
		memory[16'ha93] <= 8'hf8;
		memory[16'ha94] <= 8'h1b;
		memory[16'ha95] <= 8'h4b;
		memory[16'ha96] <= 8'h4a;
		memory[16'ha97] <= 8'h3c;
		memory[16'ha98] <= 8'h63;
		memory[16'ha99] <= 8'he7;
		memory[16'ha9a] <= 8'hdf;
		memory[16'ha9b] <= 8'h3d;
		memory[16'ha9c] <= 8'h39;
		memory[16'ha9d] <= 8'h72;
		memory[16'ha9e] <= 8'h34;
		memory[16'ha9f] <= 8'hd3;
		memory[16'haa0] <= 8'h84;
		memory[16'haa1] <= 8'he8;
		memory[16'haa2] <= 8'h80;
		memory[16'haa3] <= 8'h46;
		memory[16'haa4] <= 8'hfd;
		memory[16'haa5] <= 8'he1;
		memory[16'haa6] <= 8'h55;
		memory[16'haa7] <= 8'h27;
		memory[16'haa8] <= 8'hf;
		memory[16'haa9] <= 8'h33;
		memory[16'haaa] <= 8'h95;
		memory[16'haab] <= 8'h4a;
		memory[16'haac] <= 8'h3;
		memory[16'haad] <= 8'h17;
		memory[16'haae] <= 8'h89;
		memory[16'haaf] <= 8'hee;
		memory[16'hab0] <= 8'hf6;
		memory[16'hab1] <= 8'h72;
		memory[16'hab2] <= 8'he6;
		memory[16'hab3] <= 8'h11;
		memory[16'hab4] <= 8'hbd;
		memory[16'hab5] <= 8'h31;
		memory[16'hab6] <= 8'h4d;
		memory[16'hab7] <= 8'h20;
		memory[16'hab8] <= 8'h18;
		memory[16'hab9] <= 8'h2d;
		memory[16'haba] <= 8'h5e;
		memory[16'habb] <= 8'h52;
		memory[16'habc] <= 8'h9f;
		memory[16'habd] <= 8'h92;
		memory[16'habe] <= 8'h25;
		memory[16'habf] <= 8'h23;
		memory[16'hac0] <= 8'h7a;
		memory[16'hac1] <= 8'ha5;
		memory[16'hac2] <= 8'h69;
		memory[16'hac3] <= 8'h77;
		memory[16'hac4] <= 8'h86;
		memory[16'hac5] <= 8'hbe;
		memory[16'hac6] <= 8'h9f;
		memory[16'hac7] <= 8'h96;
		memory[16'hac8] <= 8'hf1;
		memory[16'hac9] <= 8'h34;
		memory[16'haca] <= 8'he0;
		memory[16'hacb] <= 8'hf5;
		memory[16'hacc] <= 8'h4c;
		memory[16'hacd] <= 8'h6a;
		memory[16'hace] <= 8'he3;
		memory[16'hacf] <= 8'h42;
		memory[16'had0] <= 8'hdc;
		memory[16'had1] <= 8'hca;
		memory[16'had2] <= 8'h53;
		memory[16'had3] <= 8'h9a;
		memory[16'had4] <= 8'hfb;
		memory[16'had5] <= 8'ha1;
		memory[16'had6] <= 8'hba;
		memory[16'had7] <= 8'h13;
		memory[16'had8] <= 8'hce;
		memory[16'had9] <= 8'h18;
		memory[16'hada] <= 8'h65;
		memory[16'hadb] <= 8'h6d;
		memory[16'hadc] <= 8'haa;
		memory[16'hadd] <= 8'h8a;
		memory[16'hade] <= 8'h90;
		memory[16'hadf] <= 8'h25;
		memory[16'hae0] <= 8'h30;
		memory[16'hae1] <= 8'hf9;
		memory[16'hae2] <= 8'h9c;
		memory[16'hae3] <= 8'hb6;
		memory[16'hae4] <= 8'hb8;
		memory[16'hae5] <= 8'h3b;
		memory[16'hae6] <= 8'h4c;
		memory[16'hae7] <= 8'ha9;
		memory[16'hae8] <= 8'h70;
		memory[16'hae9] <= 8'h2d;
		memory[16'haea] <= 8'h9e;
		memory[16'haeb] <= 8'hbc;
		memory[16'haec] <= 8'h97;
		memory[16'haed] <= 8'h82;
		memory[16'haee] <= 8'hfe;
		memory[16'haef] <= 8'h73;
		memory[16'haf0] <= 8'h4c;
		memory[16'haf1] <= 8'h51;
		memory[16'haf2] <= 8'hd;
		memory[16'haf3] <= 8'h47;
		memory[16'haf4] <= 8'hf2;
		memory[16'haf5] <= 8'hc8;
		memory[16'haf6] <= 8'h5a;
		memory[16'haf7] <= 8'hc0;
		memory[16'haf8] <= 8'he0;
		memory[16'haf9] <= 8'hc0;
		memory[16'hafa] <= 8'h2d;
		memory[16'hafb] <= 8'h8b;
		memory[16'hafc] <= 8'h4a;
		memory[16'hafd] <= 8'hbd;
		memory[16'hafe] <= 8'hb0;
		memory[16'haff] <= 8'h7a;
		memory[16'hb00] <= 8'hb7;
		memory[16'hb01] <= 8'h4c;
		memory[16'hb02] <= 8'h31;
		memory[16'hb03] <= 8'h6f;
		memory[16'hb04] <= 8'h88;
		memory[16'hb05] <= 8'h7d;
		memory[16'hb06] <= 8'h18;
		memory[16'hb07] <= 8'hf8;
		memory[16'hb08] <= 8'haa;
		memory[16'hb09] <= 8'hb7;
		memory[16'hb0a] <= 8'hb4;
		memory[16'hb0b] <= 8'h41;
		memory[16'hb0c] <= 8'h39;
		memory[16'hb0d] <= 8'hb2;
		memory[16'hb0e] <= 8'hb5;
		memory[16'hb0f] <= 8'h85;
		memory[16'hb10] <= 8'h3;
		memory[16'hb11] <= 8'hc2;
		memory[16'hb12] <= 8'hcc;
		memory[16'hb13] <= 8'hf6;
		memory[16'hb14] <= 8'h8a;
		memory[16'hb15] <= 8'h26;
		memory[16'hb16] <= 8'hb6;
		memory[16'hb17] <= 8'h6b;
		memory[16'hb18] <= 8'he6;
		memory[16'hb19] <= 8'he4;
		memory[16'hb1a] <= 8'hf6;
		memory[16'hb1b] <= 8'h31;
		memory[16'hb1c] <= 8'ha1;
		memory[16'hb1d] <= 8'ha6;
		memory[16'hb1e] <= 8'hab;
		memory[16'hb1f] <= 8'h58;
		memory[16'hb20] <= 8'hf2;
		memory[16'hb21] <= 8'hdc;
		memory[16'hb22] <= 8'hc7;
		memory[16'hb23] <= 8'h7a;
		memory[16'hb24] <= 8'h5a;
		memory[16'hb25] <= 8'he0;
		memory[16'hb26] <= 8'h72;
		memory[16'hb27] <= 8'h4;
		memory[16'hb28] <= 8'h97;
		memory[16'hb29] <= 8'h26;
		memory[16'hb2a] <= 8'h46;
		memory[16'hb2b] <= 8'hd0;
		memory[16'hb2c] <= 8'hd8;
		memory[16'hb2d] <= 8'hfb;
		memory[16'hb2e] <= 8'h55;
		memory[16'hb2f] <= 8'hdc;
		memory[16'hb30] <= 8'hbd;
		memory[16'hb31] <= 8'h21;
		memory[16'hb32] <= 8'hd2;
		memory[16'hb33] <= 8'h48;
		memory[16'hb34] <= 8'h47;
		memory[16'hb35] <= 8'h88;
		memory[16'hb36] <= 8'hb3;
		memory[16'hb37] <= 8'h2e;
		memory[16'hb38] <= 8'h6c;
		memory[16'hb39] <= 8'ha9;
		memory[16'hb3a] <= 8'h5f;
		memory[16'hb3b] <= 8'he;
		memory[16'hb3c] <= 8'h4f;
		memory[16'hb3d] <= 8'ha;
		memory[16'hb3e] <= 8'h66;
		memory[16'hb3f] <= 8'h41;
		memory[16'hb40] <= 8'he7;
		memory[16'hb41] <= 8'h2e;
		memory[16'hb42] <= 8'hbc;
		memory[16'hb43] <= 8'h41;
		memory[16'hb44] <= 8'he;
		memory[16'hb45] <= 8'h2e;
		memory[16'hb46] <= 8'h45;
		memory[16'hb47] <= 8'ha5;
		memory[16'hb48] <= 8'h55;
		memory[16'hb49] <= 8'h8b;
		memory[16'hb4a] <= 8'h75;
		memory[16'hb4b] <= 8'h2d;
		memory[16'hb4c] <= 8'h86;
		memory[16'hb4d] <= 8'hca;
		memory[16'hb4e] <= 8'h9;
		memory[16'hb4f] <= 8'h44;
		memory[16'hb50] <= 8'heb;
		memory[16'hb51] <= 8'hdb;
		memory[16'hb52] <= 8'h8c;
		memory[16'hb53] <= 8'h32;
		memory[16'hb54] <= 8'h64;
		memory[16'hb55] <= 8'h3f;
		memory[16'hb56] <= 8'h60;
		memory[16'hb57] <= 8'hd0;
		memory[16'hb58] <= 8'he8;
		memory[16'hb59] <= 8'hbf;
		memory[16'hb5a] <= 8'hde;
		memory[16'hb5b] <= 8'h37;
		memory[16'hb5c] <= 8'hca;
		memory[16'hb5d] <= 8'h45;
		memory[16'hb5e] <= 8'h78;
		memory[16'hb5f] <= 8'hb1;
		memory[16'hb60] <= 8'h73;
		memory[16'hb61] <= 8'h34;
		memory[16'hb62] <= 8'hf2;
		memory[16'hb63] <= 8'h81;
		memory[16'hb64] <= 8'h63;
		memory[16'hb65] <= 8'h37;
		memory[16'hb66] <= 8'h26;
		memory[16'hb67] <= 8'hb8;
		memory[16'hb68] <= 8'hc3;
		memory[16'hb69] <= 8'h9b;
		memory[16'hb6a] <= 8'he5;
		memory[16'hb6b] <= 8'h49;
		memory[16'hb6c] <= 8'h65;
		memory[16'hb6d] <= 8'hef;
		memory[16'hb6e] <= 8'h8d;
		memory[16'hb6f] <= 8'h50;
		memory[16'hb70] <= 8'hca;
		memory[16'hb71] <= 8'h19;
		memory[16'hb72] <= 8'h82;
		memory[16'hb73] <= 8'h2e;
		memory[16'hb74] <= 8'h58;
		memory[16'hb75] <= 8'he3;
		memory[16'hb76] <= 8'hff;
		memory[16'hb77] <= 8'h40;
		memory[16'hb78] <= 8'ha2;
		memory[16'hb79] <= 8'hdd;
		memory[16'hb7a] <= 8'h77;
		memory[16'hb7b] <= 8'h6c;
		memory[16'hb7c] <= 8'h22;
		memory[16'hb7d] <= 8'hf0;
		memory[16'hb7e] <= 8'h1d;
		memory[16'hb7f] <= 8'h95;
		memory[16'hb80] <= 8'h24;
		memory[16'hb81] <= 8'hf;
		memory[16'hb82] <= 8'h16;
		memory[16'hb83] <= 8'h87;
		memory[16'hb84] <= 8'h47;
		memory[16'hb85] <= 8'h3c;
		memory[16'hb86] <= 8'h3f;
		memory[16'hb87] <= 8'ha;
		memory[16'hb88] <= 8'hd7;
		memory[16'hb89] <= 8'h25;
		memory[16'hb8a] <= 8'h53;
		memory[16'hb8b] <= 8'h3c;
		memory[16'hb8c] <= 8'h14;
		memory[16'hb8d] <= 8'he1;
		memory[16'hb8e] <= 8'h8c;
		memory[16'hb8f] <= 8'hde;
		memory[16'hb90] <= 8'hfa;
		memory[16'hb91] <= 8'hf;
		memory[16'hb92] <= 8'hd;
		memory[16'hb93] <= 8'h53;
		memory[16'hb94] <= 8'hf2;
		memory[16'hb95] <= 8'hc;
		memory[16'hb96] <= 8'h93;
		memory[16'hb97] <= 8'h94;
		memory[16'hb98] <= 8'he9;
		memory[16'hb99] <= 8'hb;
		memory[16'hb9a] <= 8'h1;
		memory[16'hb9b] <= 8'hc;
		memory[16'hb9c] <= 8'hfb;
		memory[16'hb9d] <= 8'h1e;
		memory[16'hb9e] <= 8'ha1;
		memory[16'hb9f] <= 8'h1f;
		memory[16'hba0] <= 8'h2e;
		memory[16'hba1] <= 8'hb8;
		memory[16'hba2] <= 8'ha7;
		memory[16'hba3] <= 8'h75;
		memory[16'hba4] <= 8'hf4;
		memory[16'hba5] <= 8'he6;
		memory[16'hba6] <= 8'h7f;
		memory[16'hba7] <= 8'hcc;
		memory[16'hba8] <= 8'hb;
		memory[16'hba9] <= 8'hd2;
		memory[16'hbaa] <= 8'h8;
		memory[16'hbab] <= 8'h1f;
		memory[16'hbac] <= 8'hb3;
		memory[16'hbad] <= 8'h95;
		memory[16'hbae] <= 8'hfe;
		memory[16'hbaf] <= 8'hae;
		memory[16'hbb0] <= 8'ha4;
		memory[16'hbb1] <= 8'hb;
		memory[16'hbb2] <= 8'h1;
		memory[16'hbb3] <= 8'h96;
		memory[16'hbb4] <= 8'h17;
		memory[16'hbb5] <= 8'h94;
		memory[16'hbb6] <= 8'h2a;
		memory[16'hbb7] <= 8'h0;
		memory[16'hbb8] <= 8'h9f;
		memory[16'hbb9] <= 8'h2b;
		memory[16'hbba] <= 8'hc;
		memory[16'hbbb] <= 8'h9a;
		memory[16'hbbc] <= 8'h4a;
		memory[16'hbbd] <= 8'hae;
		memory[16'hbbe] <= 8'hba;
		memory[16'hbbf] <= 8'h78;
		memory[16'hbc0] <= 8'h66;
		memory[16'hbc1] <= 8'h61;
		memory[16'hbc2] <= 8'hed;
		memory[16'hbc3] <= 8'h5a;
		memory[16'hbc4] <= 8'h47;
		memory[16'hbc5] <= 8'h6c;
		memory[16'hbc6] <= 8'h26;
		memory[16'hbc7] <= 8'h53;
		memory[16'hbc8] <= 8'h3e;
		memory[16'hbc9] <= 8'h2f;
		memory[16'hbca] <= 8'h72;
		memory[16'hbcb] <= 8'hf2;
		memory[16'hbcc] <= 8'hc4;
		memory[16'hbcd] <= 8'h70;
		memory[16'hbce] <= 8'ha0;
		memory[16'hbcf] <= 8'h68;
		memory[16'hbd0] <= 8'h7b;
		memory[16'hbd1] <= 8'ha1;
		memory[16'hbd2] <= 8'hfe;
		memory[16'hbd3] <= 8'h92;
		memory[16'hbd4] <= 8'h35;
		memory[16'hbd5] <= 8'h28;
		memory[16'hbd6] <= 8'h93;
		memory[16'hbd7] <= 8'hd5;
		memory[16'hbd8] <= 8'h54;
		memory[16'hbd9] <= 8'h9f;
		memory[16'hbda] <= 8'h6f;
		memory[16'hbdb] <= 8'h9e;
		memory[16'hbdc] <= 8'h4d;
		memory[16'hbdd] <= 8'h29;
		memory[16'hbde] <= 8'h16;
		memory[16'hbdf] <= 8'hb3;
		memory[16'hbe0] <= 8'h8a;
		memory[16'hbe1] <= 8'h3;
		memory[16'hbe2] <= 8'he;
		memory[16'hbe3] <= 8'hd2;
		memory[16'hbe4] <= 8'h6f;
		memory[16'hbe5] <= 8'h34;
		memory[16'hbe6] <= 8'h25;
		memory[16'hbe7] <= 8'had;
		memory[16'hbe8] <= 8'h63;
		memory[16'hbe9] <= 8'h97;
		memory[16'hbea] <= 8'h9f;
		memory[16'hbeb] <= 8'h27;
		memory[16'hbec] <= 8'h8;
		memory[16'hbed] <= 8'h3f;
		memory[16'hbee] <= 8'h8f;
		memory[16'hbef] <= 8'h83;
		memory[16'hbf0] <= 8'he0;
		memory[16'hbf1] <= 8'h8d;
		memory[16'hbf2] <= 8'h16;
		memory[16'hbf3] <= 8'h16;
		memory[16'hbf4] <= 8'hb6;
		memory[16'hbf5] <= 8'ha9;
		memory[16'hbf6] <= 8'heb;
		memory[16'hbf7] <= 8'ha;
		memory[16'hbf8] <= 8'h48;
		memory[16'hbf9] <= 8'h5a;
		memory[16'hbfa] <= 8'ha8;
		memory[16'hbfb] <= 8'h96;
		memory[16'hbfc] <= 8'h84;
		memory[16'hbfd] <= 8'hbe;
		memory[16'hbfe] <= 8'h49;
		memory[16'hbff] <= 8'he;
		memory[16'hc00] <= 8'hc1;
		memory[16'hc01] <= 8'h57;
		memory[16'hc02] <= 8'he0;
		memory[16'hc03] <= 8'h30;
		memory[16'hc04] <= 8'h8c;
		memory[16'hc05] <= 8'h5;
		memory[16'hc06] <= 8'hdd;
		memory[16'hc07] <= 8'hef;
		memory[16'hc08] <= 8'h9d;
		memory[16'hc09] <= 8'h7d;
		memory[16'hc0a] <= 8'h17;
		memory[16'hc0b] <= 8'ha5;
		memory[16'hc0c] <= 8'hbc;
		memory[16'hc0d] <= 8'ha6;
		memory[16'hc0e] <= 8'h28;
		memory[16'hc0f] <= 8'h9d;
		memory[16'hc10] <= 8'h34;
		memory[16'hc11] <= 8'h3e;
		memory[16'hc12] <= 8'hb3;
		memory[16'hc13] <= 8'hea;
		memory[16'hc14] <= 8'he7;
		memory[16'hc15] <= 8'h9e;
		memory[16'hc16] <= 8'hf4;
		memory[16'hc17] <= 8'h30;
		memory[16'hc18] <= 8'hf8;
		memory[16'hc19] <= 8'h9c;
		memory[16'hc1a] <= 8'hc6;
		memory[16'hc1b] <= 8'h7c;
		memory[16'hc1c] <= 8'h5a;
		memory[16'hc1d] <= 8'hf;
		memory[16'hc1e] <= 8'h8b;
		memory[16'hc1f] <= 8'h1b;
		memory[16'hc20] <= 8'h67;
		memory[16'hc21] <= 8'h6b;
		memory[16'hc22] <= 8'h4b;
		memory[16'hc23] <= 8'hf3;
		memory[16'hc24] <= 8'h71;
		memory[16'hc25] <= 8'h28;
		memory[16'hc26] <= 8'he2;
		memory[16'hc27] <= 8'he;
		memory[16'hc28] <= 8'ha5;
		memory[16'hc29] <= 8'hf9;
		memory[16'hc2a] <= 8'hb3;
		memory[16'hc2b] <= 8'h62;
		memory[16'hc2c] <= 8'ha0;
		memory[16'hc2d] <= 8'hdb;
		memory[16'hc2e] <= 8'hff;
		memory[16'hc2f] <= 8'hd4;
		memory[16'hc30] <= 8'h1a;
		memory[16'hc31] <= 8'hb2;
		memory[16'hc32] <= 8'hbe;
		memory[16'hc33] <= 8'h1;
		memory[16'hc34] <= 8'h50;
		memory[16'hc35] <= 8'hb2;
		memory[16'hc36] <= 8'h31;
		memory[16'hc37] <= 8'h48;
		memory[16'hc38] <= 8'h4e;
		memory[16'hc39] <= 8'hf7;
		memory[16'hc3a] <= 8'hc5;
		memory[16'hc3b] <= 8'ha8;
		memory[16'hc3c] <= 8'h7;
		memory[16'hc3d] <= 8'h50;
		memory[16'hc3e] <= 8'hc3;
		memory[16'hc3f] <= 8'h6e;
		memory[16'hc40] <= 8'hbb;
		memory[16'hc41] <= 8'he;
		memory[16'hc42] <= 8'h61;
		memory[16'hc43] <= 8'h2c;
		memory[16'hc44] <= 8'h36;
		memory[16'hc45] <= 8'h43;
		memory[16'hc46] <= 8'h3a;
		memory[16'hc47] <= 8'hdc;
		memory[16'hc48] <= 8'h3d;
		memory[16'hc49] <= 8'hed;
		memory[16'hc4a] <= 8'h3e;
		memory[16'hc4b] <= 8'hdd;
		memory[16'hc4c] <= 8'hc9;
		memory[16'hc4d] <= 8'h3d;
		memory[16'hc4e] <= 8'hb1;
		memory[16'hc4f] <= 8'he3;
		memory[16'hc50] <= 8'hef;
		memory[16'hc51] <= 8'h6f;
		memory[16'hc52] <= 8'he4;
		memory[16'hc53] <= 8'h3f;
		memory[16'hc54] <= 8'h21;
		memory[16'hc55] <= 8'h16;
		memory[16'hc56] <= 8'h87;
		memory[16'hc57] <= 8'h6f;
		memory[16'hc58] <= 8'hd;
		memory[16'hc59] <= 8'h4c;
		memory[16'hc5a] <= 8'h17;
		memory[16'hc5b] <= 8'h14;
		memory[16'hc5c] <= 8'h9c;
		memory[16'hc5d] <= 8'hda;
		memory[16'hc5e] <= 8'h82;
		memory[16'hc5f] <= 8'h58;
		memory[16'hc60] <= 8'he8;
		memory[16'hc61] <= 8'he3;
		memory[16'hc62] <= 8'h84;
		memory[16'hc63] <= 8'h1e;
		memory[16'hc64] <= 8'h27;
		memory[16'hc65] <= 8'hbf;
		memory[16'hc66] <= 8'hfa;
		memory[16'hc67] <= 8'h64;
		memory[16'hc68] <= 8'hac;
		memory[16'hc69] <= 8'h38;
		memory[16'hc6a] <= 8'h41;
		memory[16'hc6b] <= 8'h75;
		memory[16'hc6c] <= 8'h75;
		memory[16'hc6d] <= 8'hf2;
		memory[16'hc6e] <= 8'h58;
		memory[16'hc6f] <= 8'h64;
		memory[16'hc70] <= 8'h61;
		memory[16'hc71] <= 8'h3d;
		memory[16'hc72] <= 8'ha3;
		memory[16'hc73] <= 8'h82;
		memory[16'hc74] <= 8'h53;
		memory[16'hc75] <= 8'h2b;
		memory[16'hc76] <= 8'hf1;
		memory[16'hc77] <= 8'h60;
		memory[16'hc78] <= 8'h77;
		memory[16'hc79] <= 8'h8;
		memory[16'hc7a] <= 8'h75;
		memory[16'hc7b] <= 8'h14;
		memory[16'hc7c] <= 8'he2;
		memory[16'hc7d] <= 8'hf7;
		memory[16'hc7e] <= 8'h6c;
		memory[16'hc7f] <= 8'hca;
		memory[16'hc80] <= 8'hdb;
		memory[16'hc81] <= 8'hf0;
		memory[16'hc82] <= 8'he8;
		memory[16'hc83] <= 8'h2;
		memory[16'hc84] <= 8'haf;
		memory[16'hc85] <= 8'he3;
		memory[16'hc86] <= 8'h66;
		memory[16'hc87] <= 8'h5c;
		memory[16'hc88] <= 8'h1b;
		memory[16'hc89] <= 8'ha7;
		memory[16'hc8a] <= 8'hd1;
		memory[16'hc8b] <= 8'h91;
		memory[16'hc8c] <= 8'h99;
		memory[16'hc8d] <= 8'h2a;
		memory[16'hc8e] <= 8'hf5;
		memory[16'hc8f] <= 8'hfa;
		memory[16'hc90] <= 8'h67;
		memory[16'hc91] <= 8'h99;
		memory[16'hc92] <= 8'h7c;
		memory[16'hc93] <= 8'hba;
		memory[16'hc94] <= 8'hc4;
		memory[16'hc95] <= 8'h6d;
		memory[16'hc96] <= 8'h1a;
		memory[16'hc97] <= 8'h3b;
		memory[16'hc98] <= 8'h75;
		memory[16'hc99] <= 8'h8f;
		memory[16'hc9a] <= 8'h4f;
		memory[16'hc9b] <= 8'h57;
		memory[16'hc9c] <= 8'h87;
		memory[16'hc9d] <= 8'hbb;
		memory[16'hc9e] <= 8'h21;
		memory[16'hc9f] <= 8'h62;
		memory[16'hca0] <= 8'hac;
		memory[16'hca1] <= 8'h9;
		memory[16'hca2] <= 8'h64;
		memory[16'hca3] <= 8'h5b;
		memory[16'hca4] <= 8'hec;
		memory[16'hca5] <= 8'hca;
		memory[16'hca6] <= 8'hb7;
		memory[16'hca7] <= 8'h8;
		memory[16'hca8] <= 8'h71;
		memory[16'hca9] <= 8'h89;
		memory[16'hcaa] <= 8'h99;
		memory[16'hcab] <= 8'ha;
		memory[16'hcac] <= 8'hb3;
		memory[16'hcad] <= 8'h8e;
		memory[16'hcae] <= 8'h4;
		memory[16'hcaf] <= 8'h1a;
		memory[16'hcb0] <= 8'h27;
		memory[16'hcb1] <= 8'h80;
		memory[16'hcb2] <= 8'hd4;
		memory[16'hcb3] <= 8'heb;
		memory[16'hcb4] <= 8'hed;
		memory[16'hcb5] <= 8'hee;
		memory[16'hcb6] <= 8'h27;
		memory[16'hcb7] <= 8'h62;
		memory[16'hcb8] <= 8'h7e;
		memory[16'hcb9] <= 8'h76;
		memory[16'hcba] <= 8'hb9;
		memory[16'hcbb] <= 8'h5;
		memory[16'hcbc] <= 8'h32;
		memory[16'hcbd] <= 8'hda;
		memory[16'hcbe] <= 8'h67;
		memory[16'hcbf] <= 8'hde;
		memory[16'hcc0] <= 8'he3;
		memory[16'hcc1] <= 8'hcb;
		memory[16'hcc2] <= 8'h39;
		memory[16'hcc3] <= 8'hd0;
		memory[16'hcc4] <= 8'h95;
		memory[16'hcc5] <= 8'hf1;
		memory[16'hcc6] <= 8'hd8;
		memory[16'hcc7] <= 8'h6;
		memory[16'hcc8] <= 8'h7a;
		memory[16'hcc9] <= 8'h71;
		memory[16'hcca] <= 8'h10;
		memory[16'hccb] <= 8'h2d;
		memory[16'hccc] <= 8'hff;
		memory[16'hccd] <= 8'h14;
		memory[16'hcce] <= 8'h47;
		memory[16'hccf] <= 8'h27;
		memory[16'hcd0] <= 8'h94;
		memory[16'hcd1] <= 8'h1b;
		memory[16'hcd2] <= 8'h12;
		memory[16'hcd3] <= 8'h81;
		memory[16'hcd4] <= 8'h9;
		memory[16'hcd5] <= 8'h39;
		memory[16'hcd6] <= 8'he3;
		memory[16'hcd7] <= 8'h87;
		memory[16'hcd8] <= 8'hb0;
		memory[16'hcd9] <= 8'h9c;
		memory[16'hcda] <= 8'h8c;
		memory[16'hcdb] <= 8'he2;
		memory[16'hcdc] <= 8'h76;
		memory[16'hcdd] <= 8'hf3;
		memory[16'hcde] <= 8'hc0;
		memory[16'hcdf] <= 8'h59;
		memory[16'hce0] <= 8'hbe;
		memory[16'hce1] <= 8'hf9;
		memory[16'hce2] <= 8'h29;
		memory[16'hce3] <= 8'h53;
		memory[16'hce4] <= 8'hea;
		memory[16'hce5] <= 8'h1;
		memory[16'hce6] <= 8'h59;
		memory[16'hce7] <= 8'h64;
		memory[16'hce8] <= 8'h72;
		memory[16'hce9] <= 8'h69;
		memory[16'hcea] <= 8'h91;
		memory[16'hceb] <= 8'h72;
		memory[16'hcec] <= 8'h7d;
		memory[16'hced] <= 8'hd8;
		memory[16'hcee] <= 8'h99;
		memory[16'hcef] <= 8'h11;
		memory[16'hcf0] <= 8'hf3;
		memory[16'hcf1] <= 8'hab;
		memory[16'hcf2] <= 8'h92;
		memory[16'hcf3] <= 8'hfd;
		memory[16'hcf4] <= 8'he5;
		memory[16'hcf5] <= 8'h75;
		memory[16'hcf6] <= 8'h84;
		memory[16'hcf7] <= 8'h95;
		memory[16'hcf8] <= 8'h11;
		memory[16'hcf9] <= 8'h11;
		memory[16'hcfa] <= 8'h77;
		memory[16'hcfb] <= 8'h87;
		memory[16'hcfc] <= 8'h4;
		memory[16'hcfd] <= 8'h37;
		memory[16'hcfe] <= 8'he1;
		memory[16'hcff] <= 8'hc3;
		memory[16'hd00] <= 8'h30;
		memory[16'hd01] <= 8'ha;
		memory[16'hd02] <= 8'h16;
		memory[16'hd03] <= 8'h1b;
		memory[16'hd04] <= 8'hc;
		memory[16'hd05] <= 8'h70;
		memory[16'hd06] <= 8'h7f;
		memory[16'hd07] <= 8'h7e;
		memory[16'hd08] <= 8'hd9;
		memory[16'hd09] <= 8'h11;
		memory[16'hd0a] <= 8'hf0;
		memory[16'hd0b] <= 8'h57;
		memory[16'hd0c] <= 8'he9;
		memory[16'hd0d] <= 8'h89;
		memory[16'hd0e] <= 8'h68;
		memory[16'hd0f] <= 8'hdd;
		memory[16'hd10] <= 8'h35;
		memory[16'hd11] <= 8'hfb;
		memory[16'hd12] <= 8'hda;
		memory[16'hd13] <= 8'h1a;
		memory[16'hd14] <= 8'h70;
		memory[16'hd15] <= 8'h5e;
		memory[16'hd16] <= 8'haf;
		memory[16'hd17] <= 8'h82;
		memory[16'hd18] <= 8'h6f;
		memory[16'hd19] <= 8'h26;
		memory[16'hd1a] <= 8'h9;
		memory[16'hd1b] <= 8'h74;
		memory[16'hd1c] <= 8'h5d;
		memory[16'hd1d] <= 8'hea;
		memory[16'hd1e] <= 8'h37;
		memory[16'hd1f] <= 8'h8d;
		memory[16'hd20] <= 8'hf5;
		memory[16'hd21] <= 8'h4d;
		memory[16'hd22] <= 8'ha8;
		memory[16'hd23] <= 8'h1;
		memory[16'hd24] <= 8'hbd;
		memory[16'hd25] <= 8'h28;
		memory[16'hd26] <= 8'h7f;
		memory[16'hd27] <= 8'h97;
		memory[16'hd28] <= 8'h39;
		memory[16'hd29] <= 8'h70;
		memory[16'hd2a] <= 8'hee;
		memory[16'hd2b] <= 8'h22;
		memory[16'hd2c] <= 8'hf9;
		memory[16'hd2d] <= 8'h56;
		memory[16'hd2e] <= 8'hff;
		memory[16'hd2f] <= 8'h2e;
		memory[16'hd30] <= 8'h51;
		memory[16'hd31] <= 8'hd9;
		memory[16'hd32] <= 8'h48;
		memory[16'hd33] <= 8'hc2;
		memory[16'hd34] <= 8'h38;
		memory[16'hd35] <= 8'hf7;
		memory[16'hd36] <= 8'h44;
		memory[16'hd37] <= 8'ha7;
		memory[16'hd38] <= 8'h1d;
		memory[16'hd39] <= 8'h4d;
		memory[16'hd3a] <= 8'h1b;
		memory[16'hd3b] <= 8'h7a;
		memory[16'hd3c] <= 8'h38;
		memory[16'hd3d] <= 8'h52;
		memory[16'hd3e] <= 8'h8;
		memory[16'hd3f] <= 8'h2d;
		memory[16'hd40] <= 8'ha0;
		memory[16'hd41] <= 8'hb0;
		memory[16'hd42] <= 8'h2e;
		memory[16'hd43] <= 8'h5d;
		memory[16'hd44] <= 8'hd8;
		memory[16'hd45] <= 8'had;
		memory[16'hd46] <= 8'hf4;
		memory[16'hd47] <= 8'h11;
		memory[16'hd48] <= 8'h1d;
		memory[16'hd49] <= 8'he2;
		memory[16'hd4a] <= 8'h34;
		memory[16'hd4b] <= 8'h17;
		memory[16'hd4c] <= 8'h39;
		memory[16'hd4d] <= 8'h33;
		memory[16'hd4e] <= 8'h45;
		memory[16'hd4f] <= 8'h8a;
		memory[16'hd50] <= 8'hd;
		memory[16'hd51] <= 8'h8e;
		memory[16'hd52] <= 8'h4c;
		memory[16'hd53] <= 8'h45;
		memory[16'hd54] <= 8'h85;
		memory[16'hd55] <= 8'h90;
		memory[16'hd56] <= 8'hec;
		memory[16'hd57] <= 8'ha3;
		memory[16'hd58] <= 8'hde;
		memory[16'hd59] <= 8'h8;
		memory[16'hd5a] <= 8'h1d;
		memory[16'hd5b] <= 8'h16;
		memory[16'hd5c] <= 8'h5a;
		memory[16'hd5d] <= 8'h25;
		memory[16'hd5e] <= 8'h43;
		memory[16'hd5f] <= 8'hfa;
		memory[16'hd60] <= 8'hd6;
		memory[16'hd61] <= 8'h71;
		memory[16'hd62] <= 8'h58;
		memory[16'hd63] <= 8'hae;
		memory[16'hd64] <= 8'h1e;
		memory[16'hd65] <= 8'h4c;
		memory[16'hd66] <= 8'hc0;
		memory[16'hd67] <= 8'h3c;
		memory[16'hd68] <= 8'h2f;
		memory[16'hd69] <= 8'hf4;
		memory[16'hd6a] <= 8'h53;
		memory[16'hd6b] <= 8'h68;
		memory[16'hd6c] <= 8'h27;
		memory[16'hd6d] <= 8'h98;
		memory[16'hd6e] <= 8'hf2;
		memory[16'hd6f] <= 8'h34;
		memory[16'hd70] <= 8'h26;
		memory[16'hd71] <= 8'h3f;
		memory[16'hd72] <= 8'h79;
		memory[16'hd73] <= 8'hac;
		memory[16'hd74] <= 8'hcf;
		memory[16'hd75] <= 8'h66;
		memory[16'hd76] <= 8'h4f;
		memory[16'hd77] <= 8'had;
		memory[16'hd78] <= 8'h6e;
		memory[16'hd79] <= 8'h6c;
		memory[16'hd7a] <= 8'hc3;
		memory[16'hd7b] <= 8'hc8;
		memory[16'hd7c] <= 8'h92;
		memory[16'hd7d] <= 8'h6;
		memory[16'hd7e] <= 8'hc3;
		memory[16'hd7f] <= 8'h68;
		memory[16'hd80] <= 8'h77;
		memory[16'hd81] <= 8'h1b;
		memory[16'hd82] <= 8'h16;
		memory[16'hd83] <= 8'h96;
		memory[16'hd84] <= 8'h67;
		memory[16'hd85] <= 8'hd6;
		memory[16'hd86] <= 8'hd2;
		memory[16'hd87] <= 8'h96;
		memory[16'hd88] <= 8'hca;
		memory[16'hd89] <= 8'h25;
		memory[16'hd8a] <= 8'hfe;
		memory[16'hd8b] <= 8'hf2;
		memory[16'hd8c] <= 8'hbd;
		memory[16'hd8d] <= 8'hf1;
		memory[16'hd8e] <= 8'h26;
		memory[16'hd8f] <= 8'he4;
		memory[16'hd90] <= 8'h30;
		memory[16'hd91] <= 8'ha0;
		memory[16'hd92] <= 8'h90;
		memory[16'hd93] <= 8'hff;
		memory[16'hd94] <= 8'h6;
		memory[16'hd95] <= 8'hdf;
		memory[16'hd96] <= 8'had;
		memory[16'hd97] <= 8'h74;
		memory[16'hd98] <= 8'h4b;
		memory[16'hd99] <= 8'h70;
		memory[16'hd9a] <= 8'h3c;
		memory[16'hd9b] <= 8'hdd;
		memory[16'hd9c] <= 8'h77;
		memory[16'hd9d] <= 8'hff;
		memory[16'hd9e] <= 8'h45;
		memory[16'hd9f] <= 8'hee;
		memory[16'hda0] <= 8'h1a;
		memory[16'hda1] <= 8'h5c;
		memory[16'hda2] <= 8'h84;
		memory[16'hda3] <= 8'h82;
		memory[16'hda4] <= 8'h32;
		memory[16'hda5] <= 8'h56;
		memory[16'hda6] <= 8'h18;
		memory[16'hda7] <= 8'hfd;
		memory[16'hda8] <= 8'h7b;
		memory[16'hda9] <= 8'h17;
		memory[16'hdaa] <= 8'hef;
		memory[16'hdab] <= 8'h39;
		memory[16'hdac] <= 8'h8;
		memory[16'hdad] <= 8'h15;
		memory[16'hdae] <= 8'h1d;
		memory[16'hdaf] <= 8'h38;
		memory[16'hdb0] <= 8'hb5;
		memory[16'hdb1] <= 8'had;
		memory[16'hdb2] <= 8'h37;
		memory[16'hdb3] <= 8'hbb;
		memory[16'hdb4] <= 8'h8c;
		memory[16'hdb5] <= 8'he4;
		memory[16'hdb6] <= 8'h2f;
		memory[16'hdb7] <= 8'hd7;
		memory[16'hdb8] <= 8'h55;
		memory[16'hdb9] <= 8'h6c;
		memory[16'hdba] <= 8'hb5;
		memory[16'hdbb] <= 8'hcc;
		memory[16'hdbc] <= 8'h6b;
		memory[16'hdbd] <= 8'hfa;
		memory[16'hdbe] <= 8'hba;
		memory[16'hdbf] <= 8'h86;
		memory[16'hdc0] <= 8'h56;
		memory[16'hdc1] <= 8'h3f;
		memory[16'hdc2] <= 8'h8;
		memory[16'hdc3] <= 8'h89;
		memory[16'hdc4] <= 8'h95;
		memory[16'hdc5] <= 8'h20;
		memory[16'hdc6] <= 8'h86;
		memory[16'hdc7] <= 8'h11;
		memory[16'hdc8] <= 8'h37;
		memory[16'hdc9] <= 8'h75;
		memory[16'hdca] <= 8'h4a;
		memory[16'hdcb] <= 8'h3f;
		memory[16'hdcc] <= 8'h8a;
		memory[16'hdcd] <= 8'h67;
		memory[16'hdce] <= 8'h77;
		memory[16'hdcf] <= 8'h40;
		memory[16'hdd0] <= 8'h14;
		memory[16'hdd1] <= 8'haf;
		memory[16'hdd2] <= 8'hfb;
		memory[16'hdd3] <= 8'ha0;
		memory[16'hdd4] <= 8'h93;
		memory[16'hdd5] <= 8'h2b;
		memory[16'hdd6] <= 8'h77;
		memory[16'hdd7] <= 8'he8;
		memory[16'hdd8] <= 8'h97;
		memory[16'hdd9] <= 8'h2c;
		memory[16'hdda] <= 8'hb4;
		memory[16'hddb] <= 8'h2;
		memory[16'hddc] <= 8'h27;
		memory[16'hddd] <= 8'h6f;
		memory[16'hdde] <= 8'h88;
		memory[16'hddf] <= 8'h7d;
		memory[16'hde0] <= 8'hae;
		memory[16'hde1] <= 8'h90;
		memory[16'hde2] <= 8'h6;
		memory[16'hde3] <= 8'h43;
		memory[16'hde4] <= 8'hb1;
		memory[16'hde5] <= 8'h8c;
		memory[16'hde6] <= 8'h54;
		memory[16'hde7] <= 8'he8;
		memory[16'hde8] <= 8'h1;
		memory[16'hde9] <= 8'h9e;
		memory[16'hdea] <= 8'h28;
		memory[16'hdeb] <= 8'h8c;
		memory[16'hdec] <= 8'h5;
		memory[16'hded] <= 8'h9f;
		memory[16'hdee] <= 8'hcc;
		memory[16'hdef] <= 8'h19;
		memory[16'hdf0] <= 8'h4e;
		memory[16'hdf1] <= 8'hc7;
		memory[16'hdf2] <= 8'hb9;
		memory[16'hdf3] <= 8'he2;
		memory[16'hdf4] <= 8'hf2;
		memory[16'hdf5] <= 8'h31;
		memory[16'hdf6] <= 8'hca;
		memory[16'hdf7] <= 8'h89;
		memory[16'hdf8] <= 8'h5d;
		memory[16'hdf9] <= 8'h7f;
		memory[16'hdfa] <= 8'h8c;
		memory[16'hdfb] <= 8'h84;
		memory[16'hdfc] <= 8'hee;
		memory[16'hdfd] <= 8'h14;
		memory[16'hdfe] <= 8'h2;
		memory[16'hdff] <= 8'h9c;
		memory[16'he00] <= 8'ha5;
		memory[16'he01] <= 8'h8;
		memory[16'he02] <= 8'hdf;
		memory[16'he03] <= 8'h56;
		memory[16'he04] <= 8'h95;
		memory[16'he05] <= 8'h34;
		memory[16'he06] <= 8'h3e;
		memory[16'he07] <= 8'h96;
		memory[16'he08] <= 8'hd2;
		memory[16'he09] <= 8'h66;
		memory[16'he0a] <= 8'h22;
		memory[16'he0b] <= 8'hd8;
		memory[16'he0c] <= 8'h6;
		memory[16'he0d] <= 8'hee;
		memory[16'he0e] <= 8'hf1;
		memory[16'he0f] <= 8'h54;
		memory[16'he10] <= 8'hb6;
		memory[16'he11] <= 8'hab;
		memory[16'he12] <= 8'h36;
		memory[16'he13] <= 8'ha8;
		memory[16'he14] <= 8'hdc;
		memory[16'he15] <= 8'h1;
		memory[16'he16] <= 8'h32;
		memory[16'he17] <= 8'h39;
		memory[16'he18] <= 8'h80;
		memory[16'he19] <= 8'hbe;
		memory[16'he1a] <= 8'hbe;
		memory[16'he1b] <= 8'h6e;
		memory[16'he1c] <= 8'hd2;
		memory[16'he1d] <= 8'hc0;
		memory[16'he1e] <= 8'ha;
		memory[16'he1f] <= 8'h77;
		memory[16'he20] <= 8'hc8;
		memory[16'he21] <= 8'he9;
		memory[16'he22] <= 8'hcd;
		memory[16'he23] <= 8'h5d;
		memory[16'he24] <= 8'h1d;
		memory[16'he25] <= 8'hc;
		memory[16'he26] <= 8'hf4;
		memory[16'he27] <= 8'hf0;
		memory[16'he28] <= 8'h72;
		memory[16'he29] <= 8'h16;
		memory[16'he2a] <= 8'hc8;
		memory[16'he2b] <= 8'h78;
		memory[16'he2c] <= 8'h5;
		memory[16'he2d] <= 8'hb9;
		memory[16'he2e] <= 8'hcd;
		memory[16'he2f] <= 8'hbb;
		memory[16'he30] <= 8'h64;
		memory[16'he31] <= 8'h3;
		memory[16'he32] <= 8'h63;
		memory[16'he33] <= 8'h40;
		memory[16'he34] <= 8'h4;
		memory[16'he35] <= 8'h95;
		memory[16'he36] <= 8'h7a;
		memory[16'he37] <= 8'h84;
		memory[16'he38] <= 8'h53;
		memory[16'he39] <= 8'h38;
		memory[16'he3a] <= 8'hf2;
		memory[16'he3b] <= 8'h26;
		memory[16'he3c] <= 8'hf8;
		memory[16'he3d] <= 8'hfc;
		memory[16'he3e] <= 8'h9d;
		memory[16'he3f] <= 8'hc0;
		memory[16'he40] <= 8'he6;
		memory[16'he41] <= 8'h6b;
		memory[16'he42] <= 8'h1e;
		memory[16'he43] <= 8'h3;
		memory[16'he44] <= 8'h77;
		memory[16'he45] <= 8'h12;
		memory[16'he46] <= 8'hf3;
		memory[16'he47] <= 8'he9;
		memory[16'he48] <= 8'h28;
		memory[16'he49] <= 8'hbb;
		memory[16'he4a] <= 8'h62;
		memory[16'he4b] <= 8'h2d;
		memory[16'he4c] <= 8'h75;
		memory[16'he4d] <= 8'h2f;
		memory[16'he4e] <= 8'he8;
		memory[16'he4f] <= 8'hd9;
		memory[16'he50] <= 8'h32;
		memory[16'he51] <= 8'h4c;
		memory[16'he52] <= 8'h1a;
		memory[16'he53] <= 8'h37;
		memory[16'he54] <= 8'he1;
		memory[16'he55] <= 8'h94;
		memory[16'he56] <= 8'hbb;
		memory[16'he57] <= 8'h35;
		memory[16'he58] <= 8'hcc;
		memory[16'he59] <= 8'hae;
		memory[16'he5a] <= 8'h5b;
		memory[16'he5b] <= 8'hc4;
		memory[16'he5c] <= 8'haa;
		memory[16'he5d] <= 8'hf8;
		memory[16'he5e] <= 8'h84;
		memory[16'he5f] <= 8'h90;
		memory[16'he60] <= 8'h63;
		memory[16'he61] <= 8'ha2;
		memory[16'he62] <= 8'h94;
		memory[16'he63] <= 8'hda;
		memory[16'he64] <= 8'hb4;
		memory[16'he65] <= 8'h87;
		memory[16'he66] <= 8'hc4;
		memory[16'he67] <= 8'hdd;
		memory[16'he68] <= 8'h43;
		memory[16'he69] <= 8'h26;
		memory[16'he6a] <= 8'ha;
		memory[16'he6b] <= 8'hb8;
		memory[16'he6c] <= 8'h55;
		memory[16'he6d] <= 8'hf3;
		memory[16'he6e] <= 8'h91;
		memory[16'he6f] <= 8'h87;
		memory[16'he70] <= 8'h3f;
		memory[16'he71] <= 8'hab;
		memory[16'he72] <= 8'hbe;
		memory[16'he73] <= 8'h20;
		memory[16'he74] <= 8'h3f;
		memory[16'he75] <= 8'h7a;
		memory[16'he76] <= 8'h55;
		memory[16'he77] <= 8'hb;
		memory[16'he78] <= 8'h28;
		memory[16'he79] <= 8'hb0;
		memory[16'he7a] <= 8'hcf;
		memory[16'he7b] <= 8'hd2;
		memory[16'he7c] <= 8'ha9;
		memory[16'he7d] <= 8'h54;
		memory[16'he7e] <= 8'h63;
		memory[16'he7f] <= 8'hc;
		memory[16'he80] <= 8'hf6;
		memory[16'he81] <= 8'hf7;
		memory[16'he82] <= 8'he7;
		memory[16'he83] <= 8'hab;
		memory[16'he84] <= 8'h7e;
		memory[16'he85] <= 8'hab;
		memory[16'he86] <= 8'h88;
		memory[16'he87] <= 8'hc1;
		memory[16'he88] <= 8'hd1;
		memory[16'he89] <= 8'h92;
		memory[16'he8a] <= 8'h79;
		memory[16'he8b] <= 8'h26;
		memory[16'he8c] <= 8'h85;
		memory[16'he8d] <= 8'hb;
		memory[16'he8e] <= 8'had;
		memory[16'he8f] <= 8'hc4;
		memory[16'he90] <= 8'hb6;
		memory[16'he91] <= 8'h6c;
		memory[16'he92] <= 8'he5;
		memory[16'he93] <= 8'hf6;
		memory[16'he94] <= 8'he6;
		memory[16'he95] <= 8'h3a;
		memory[16'he96] <= 8'h1;
		memory[16'he97] <= 8'he;
		memory[16'he98] <= 8'heb;
		memory[16'he99] <= 8'hd1;
		memory[16'he9a] <= 8'he0;
		memory[16'he9b] <= 8'h94;
		memory[16'he9c] <= 8'h25;
		memory[16'he9d] <= 8'h43;
		memory[16'he9e] <= 8'ha0;
		memory[16'he9f] <= 8'h1b;
		memory[16'hea0] <= 8'h3a;
		memory[16'hea1] <= 8'h87;
		memory[16'hea2] <= 8'hc6;
		memory[16'hea3] <= 8'hb9;
		memory[16'hea4] <= 8'h32;
		memory[16'hea5] <= 8'h4e;
		memory[16'hea6] <= 8'h7a;
		memory[16'hea7] <= 8'h3;
		memory[16'hea8] <= 8'he1;
		memory[16'hea9] <= 8'hf4;
		memory[16'heaa] <= 8'h29;
		memory[16'heab] <= 8'h66;
		memory[16'heac] <= 8'hff;
		memory[16'head] <= 8'hd7;
		memory[16'heae] <= 8'h2b;
		memory[16'heaf] <= 8'hb5;
		memory[16'heb0] <= 8'h43;
		memory[16'heb1] <= 8'h10;
		memory[16'heb2] <= 8'hab;
		memory[16'heb3] <= 8'h29;
		memory[16'heb4] <= 8'h4a;
		memory[16'heb5] <= 8'had;
		memory[16'heb6] <= 8'h37;
		memory[16'heb7] <= 8'h35;
		memory[16'heb8] <= 8'h7e;
		memory[16'heb9] <= 8'h17;
		memory[16'heba] <= 8'hc9;
		memory[16'hebb] <= 8'ha3;
		memory[16'hebc] <= 8'h5b;
		memory[16'hebd] <= 8'h6a;
		memory[16'hebe] <= 8'hbe;
		memory[16'hebf] <= 8'h95;
		memory[16'hec0] <= 8'hf1;
		memory[16'hec1] <= 8'h85;
		memory[16'hec2] <= 8'h4e;
		memory[16'hec3] <= 8'h24;
		memory[16'hec4] <= 8'hd3;
		memory[16'hec5] <= 8'hc9;
		memory[16'hec6] <= 8'h27;
		memory[16'hec7] <= 8'hb4;
		memory[16'hec8] <= 8'hbd;
		memory[16'hec9] <= 8'h51;
		memory[16'heca] <= 8'h1b;
		memory[16'hecb] <= 8'hbc;
		memory[16'hecc] <= 8'h28;
		memory[16'hecd] <= 8'h46;
		memory[16'hece] <= 8'h71;
		memory[16'hecf] <= 8'h6b;
		memory[16'hed0] <= 8'h56;
		memory[16'hed1] <= 8'h1d;
		memory[16'hed2] <= 8'h94;
		memory[16'hed3] <= 8'ha0;
		memory[16'hed4] <= 8'hca;
		memory[16'hed5] <= 8'hcb;
		memory[16'hed6] <= 8'hd6;
		memory[16'hed7] <= 8'h48;
		memory[16'hed8] <= 8'he2;
		memory[16'hed9] <= 8'h9f;
		memory[16'heda] <= 8'heb;
		memory[16'hedb] <= 8'h3d;
		memory[16'hedc] <= 8'h9;
		memory[16'hedd] <= 8'ha9;
		memory[16'hede] <= 8'hd3;
		memory[16'hedf] <= 8'hfb;
		memory[16'hee0] <= 8'h2e;
		memory[16'hee1] <= 8'h21;
		memory[16'hee2] <= 8'h1f;
		memory[16'hee3] <= 8'h2;
		memory[16'hee4] <= 8'hea;
		memory[16'hee5] <= 8'h46;
		memory[16'hee6] <= 8'hb6;
		memory[16'hee7] <= 8'ha7;
		memory[16'hee8] <= 8'h97;
		memory[16'hee9] <= 8'hd1;
		memory[16'heea] <= 8'h63;
		memory[16'heeb] <= 8'hbf;
		memory[16'heec] <= 8'h17;
		memory[16'heed] <= 8'hd5;
		memory[16'heee] <= 8'h2a;
		memory[16'heef] <= 8'h6d;
		memory[16'hef0] <= 8'hf2;
		memory[16'hef1] <= 8'hbe;
		memory[16'hef2] <= 8'he;
		memory[16'hef3] <= 8'hbc;
		memory[16'hef4] <= 8'h89;
		memory[16'hef5] <= 8'he4;
		memory[16'hef6] <= 8'h4;
		memory[16'hef7] <= 8'h6c;
		memory[16'hef8] <= 8'h83;
		memory[16'hef9] <= 8'hef;
		memory[16'hefa] <= 8'ha9;
		memory[16'hefb] <= 8'h8d;
		memory[16'hefc] <= 8'h98;
		memory[16'hefd] <= 8'h7c;
		memory[16'hefe] <= 8'h88;
		memory[16'heff] <= 8'hc7;
		memory[16'hf00] <= 8'h9e;
		memory[16'hf01] <= 8'ha7;
		memory[16'hf02] <= 8'hc9;
		memory[16'hf03] <= 8'h88;
		memory[16'hf04] <= 8'hed;
		memory[16'hf05] <= 8'h7f;
		memory[16'hf06] <= 8'h30;
		memory[16'hf07] <= 8'h85;
		memory[16'hf08] <= 8'h51;
		memory[16'hf09] <= 8'h93;
		memory[16'hf0a] <= 8'h44;
		memory[16'hf0b] <= 8'h68;
		memory[16'hf0c] <= 8'h68;
		memory[16'hf0d] <= 8'h6f;
		memory[16'hf0e] <= 8'hd6;
		memory[16'hf0f] <= 8'h5a;
		memory[16'hf10] <= 8'h2d;
		memory[16'hf11] <= 8'he4;
		memory[16'hf12] <= 8'h16;
		memory[16'hf13] <= 8'hb7;
		memory[16'hf14] <= 8'hc8;
		memory[16'hf15] <= 8'h1a;
		memory[16'hf16] <= 8'h23;
		memory[16'hf17] <= 8'h4b;
		memory[16'hf18] <= 8'h9;
		memory[16'hf19] <= 8'hcc;
		memory[16'hf1a] <= 8'hd8;
		memory[16'hf1b] <= 8'ha2;
		memory[16'hf1c] <= 8'h49;
		memory[16'hf1d] <= 8'h60;
		memory[16'hf1e] <= 8'h69;
		memory[16'hf1f] <= 8'he7;
		memory[16'hf20] <= 8'h7;
		memory[16'hf21] <= 8'h32;
		memory[16'hf22] <= 8'h6f;
		memory[16'hf23] <= 8'hf5;
		memory[16'hf24] <= 8'hb1;
		memory[16'hf25] <= 8'h9f;
		memory[16'hf26] <= 8'h7a;
		memory[16'hf27] <= 8'h2;
		memory[16'hf28] <= 8'h33;
		memory[16'hf29] <= 8'hbe;
		memory[16'hf2a] <= 8'h6b;
		memory[16'hf2b] <= 8'h9b;
		memory[16'hf2c] <= 8'h2d;
		memory[16'hf2d] <= 8'h41;
		memory[16'hf2e] <= 8'hf6;
		memory[16'hf2f] <= 8'h5b;
		memory[16'hf30] <= 8'h25;
		memory[16'hf31] <= 8'hc;
		memory[16'hf32] <= 8'h12;
		memory[16'hf33] <= 8'hed;
		memory[16'hf34] <= 8'h27;
		memory[16'hf35] <= 8'h35;
		memory[16'hf36] <= 8'h38;
		memory[16'hf37] <= 8'h30;
		memory[16'hf38] <= 8'h1;
		memory[16'hf39] <= 8'h11;
		memory[16'hf3a] <= 8'hd2;
		memory[16'hf3b] <= 8'h4a;
		memory[16'hf3c] <= 8'h71;
		memory[16'hf3d] <= 8'h3b;
		memory[16'hf3e] <= 8'h31;
		memory[16'hf3f] <= 8'h79;
		memory[16'hf40] <= 8'h6d;
		memory[16'hf41] <= 8'ha1;
		memory[16'hf42] <= 8'h6e;
		memory[16'hf43] <= 8'h1f;
		memory[16'hf44] <= 8'h40;
		memory[16'hf45] <= 8'he8;
		memory[16'hf46] <= 8'h21;
		memory[16'hf47] <= 8'h73;
		memory[16'hf48] <= 8'ha6;
		memory[16'hf49] <= 8'h8c;
		memory[16'hf4a] <= 8'hf;
		memory[16'hf4b] <= 8'hd4;
		memory[16'hf4c] <= 8'hcd;
		memory[16'hf4d] <= 8'h5;
		memory[16'hf4e] <= 8'h2f;
		memory[16'hf4f] <= 8'hf2;
		memory[16'hf50] <= 8'h11;
		memory[16'hf51] <= 8'h41;
		memory[16'hf52] <= 8'hdf;
		memory[16'hf53] <= 8'h38;
		memory[16'hf54] <= 8'h76;
		memory[16'hf55] <= 8'h18;
		memory[16'hf56] <= 8'h69;
		memory[16'hf57] <= 8'h77;
		memory[16'hf58] <= 8'h29;
		memory[16'hf59] <= 8'h3b;
		memory[16'hf5a] <= 8'hc2;
		memory[16'hf5b] <= 8'h9a;
		memory[16'hf5c] <= 8'h77;
		memory[16'hf5d] <= 8'hf3;
		memory[16'hf5e] <= 8'h13;
		memory[16'hf5f] <= 8'he4;
		memory[16'hf60] <= 8'h94;
		memory[16'hf61] <= 8'h81;
		memory[16'hf62] <= 8'h3;
		memory[16'hf63] <= 8'hd5;
		memory[16'hf64] <= 8'h69;
		memory[16'hf65] <= 8'h25;
		memory[16'hf66] <= 8'h48;
		memory[16'hf67] <= 8'h10;
		memory[16'hf68] <= 8'hb1;
		memory[16'hf69] <= 8'h57;
		memory[16'hf6a] <= 8'he4;
		memory[16'hf6b] <= 8'h7f;
		memory[16'hf6c] <= 8'h5c;
		memory[16'hf6d] <= 8'h13;
		memory[16'hf6e] <= 8'h71;
		memory[16'hf6f] <= 8'h6e;
		memory[16'hf70] <= 8'h54;
		memory[16'hf71] <= 8'h51;
		memory[16'hf72] <= 8'ha6;
		memory[16'hf73] <= 8'hca;
		memory[16'hf74] <= 8'h69;
		memory[16'hf75] <= 8'hf;
		memory[16'hf76] <= 8'h41;
		memory[16'hf77] <= 8'h92;
		memory[16'hf78] <= 8'h4b;
		memory[16'hf79] <= 8'h3;
		memory[16'hf7a] <= 8'h2c;
		memory[16'hf7b] <= 8'hc2;
		memory[16'hf7c] <= 8'hf7;
		memory[16'hf7d] <= 8'h40;
		memory[16'hf7e] <= 8'ha6;
		memory[16'hf7f] <= 8'h8b;
		memory[16'hf80] <= 8'hc1;
		memory[16'hf81] <= 8'haa;
		memory[16'hf82] <= 8'h60;
		memory[16'hf83] <= 8'h2b;
		memory[16'hf84] <= 8'hcf;
		memory[16'hf85] <= 8'ha9;
		memory[16'hf86] <= 8'h3b;
		memory[16'hf87] <= 8'h80;
		memory[16'hf88] <= 8'h0;
		memory[16'hf89] <= 8'h1f;
		memory[16'hf8a] <= 8'hff;
		memory[16'hf8b] <= 8'h5d;
		memory[16'hf8c] <= 8'h32;
		memory[16'hf8d] <= 8'h71;
		memory[16'hf8e] <= 8'hcb;
		memory[16'hf8f] <= 8'h86;
		memory[16'hf90] <= 8'hc2;
		memory[16'hf91] <= 8'h71;
		memory[16'hf92] <= 8'h50;
		memory[16'hf93] <= 8'h2b;
		memory[16'hf94] <= 8'h81;
		memory[16'hf95] <= 8'h91;
		memory[16'hf96] <= 8'hbd;
		memory[16'hf97] <= 8'hcc;
		memory[16'hf98] <= 8'h95;
		memory[16'hf99] <= 8'he9;
		memory[16'hf9a] <= 8'h8e;
		memory[16'hf9b] <= 8'h8c;
		memory[16'hf9c] <= 8'h29;
		memory[16'hf9d] <= 8'h34;
		memory[16'hf9e] <= 8'h17;
		memory[16'hf9f] <= 8'heb;
		memory[16'hfa0] <= 8'hde;
		memory[16'hfa1] <= 8'h78;
		memory[16'hfa2] <= 8'h16;
		memory[16'hfa3] <= 8'had;
		memory[16'hfa4] <= 8'h21;
		memory[16'hfa5] <= 8'h51;
		memory[16'hfa6] <= 8'h2e;
		memory[16'hfa7] <= 8'h21;
		memory[16'hfa8] <= 8'h70;
		memory[16'hfa9] <= 8'h2d;
		memory[16'hfaa] <= 8'h7e;
		memory[16'hfab] <= 8'ha2;
		memory[16'hfac] <= 8'h9e;
		memory[16'hfad] <= 8'h49;
		memory[16'hfae] <= 8'h28;
		memory[16'hfaf] <= 8'h60;
		memory[16'hfb0] <= 8'hbb;
		memory[16'hfb1] <= 8'h78;
		memory[16'hfb2] <= 8'h8b;
		memory[16'hfb3] <= 8'h3c;
		memory[16'hfb4] <= 8'h9;
		memory[16'hfb5] <= 8'h48;
		memory[16'hfb6] <= 8'h8;
		memory[16'hfb7] <= 8'h9e;
		memory[16'hfb8] <= 8'h32;
		memory[16'hfb9] <= 8'h96;
		memory[16'hfba] <= 8'h2a;
		memory[16'hfbb] <= 8'h5b;
		memory[16'hfbc] <= 8'hca;
		memory[16'hfbd] <= 8'h42;
		memory[16'hfbe] <= 8'h46;
		memory[16'hfbf] <= 8'ha9;
		memory[16'hfc0] <= 8'hba;
		memory[16'hfc1] <= 8'h5c;
		memory[16'hfc2] <= 8'h56;
		memory[16'hfc3] <= 8'hdb;
		memory[16'hfc4] <= 8'had;
		memory[16'hfc5] <= 8'h84;
		memory[16'hfc6] <= 8'hfc;
		memory[16'hfc7] <= 8'h1d;
		memory[16'hfc8] <= 8'hb2;
		memory[16'hfc9] <= 8'h7b;
		memory[16'hfca] <= 8'hbf;
		memory[16'hfcb] <= 8'h50;
		memory[16'hfcc] <= 8'hc4;
		memory[16'hfcd] <= 8'he7;
		memory[16'hfce] <= 8'hb1;
		memory[16'hfcf] <= 8'h7f;
		memory[16'hfd0] <= 8'h5f;
		memory[16'hfd1] <= 8'h3c;
		memory[16'hfd2] <= 8'hbb;
		memory[16'hfd3] <= 8'h69;
		memory[16'hfd4] <= 8'h85;
		memory[16'hfd5] <= 8'hc3;
		memory[16'hfd6] <= 8'h7;
		memory[16'hfd7] <= 8'hb7;
		memory[16'hfd8] <= 8'h59;
		memory[16'hfd9] <= 8'h32;
		memory[16'hfda] <= 8'h12;
		memory[16'hfdb] <= 8'h24;
		memory[16'hfdc] <= 8'h74;
		memory[16'hfdd] <= 8'h59;
		memory[16'hfde] <= 8'hcd;
		memory[16'hfdf] <= 8'h2e;
		memory[16'hfe0] <= 8'hb5;
		memory[16'hfe1] <= 8'h23;
		memory[16'hfe2] <= 8'h9;
		memory[16'hfe3] <= 8'h63;
		memory[16'hfe4] <= 8'ha8;
		memory[16'hfe5] <= 8'h5;
		memory[16'hfe6] <= 8'h80;
		memory[16'hfe7] <= 8'h5a;
		memory[16'hfe8] <= 8'h80;
		memory[16'hfe9] <= 8'h40;
		memory[16'hfea] <= 8'haa;
		memory[16'hfeb] <= 8'h45;
		memory[16'hfec] <= 8'h27;
		memory[16'hfed] <= 8'h5b;
		memory[16'hfee] <= 8'hc4;
		memory[16'hfef] <= 8'h87;
		memory[16'hff0] <= 8'h98;
		memory[16'hff1] <= 8'h80;
		memory[16'hff2] <= 8'hf0;
		memory[16'hff3] <= 8'h1d;
		memory[16'hff4] <= 8'h43;
		memory[16'hff5] <= 8'hf7;
		memory[16'hff6] <= 8'hd4;
		memory[16'hff7] <= 8'h9d;
		memory[16'hff8] <= 8'h29;
		memory[16'hff9] <= 8'he6;
		memory[16'hffa] <= 8'hc1;
		memory[16'hffb] <= 8'h9d;
		memory[16'hffc] <= 8'h3f;
		memory[16'hffd] <= 8'h8e;
		memory[16'hffe] <= 8'hcb;
		memory[16'hfff] <= 8'hf5;
		memory[16'h1000] <= 8'hb1;
		memory[16'h1001] <= 8'hd4;
		memory[16'h1002] <= 8'h58;
		memory[16'h1003] <= 8'h59;
		memory[16'h1004] <= 8'hda;
		memory[16'h1005] <= 8'hd8;
		memory[16'h1006] <= 8'hb3;
		memory[16'h1007] <= 8'h5a;
		memory[16'h1008] <= 8'h18;
		memory[16'h1009] <= 8'h5e;
		memory[16'h100a] <= 8'h9f;
		memory[16'h100b] <= 8'h40;
		memory[16'h100c] <= 8'hb9;
		memory[16'h100d] <= 8'h64;
		memory[16'h100e] <= 8'hc7;
		memory[16'h100f] <= 8'h51;
		memory[16'h1010] <= 8'he4;
		memory[16'h1011] <= 8'hb7;
		memory[16'h1012] <= 8'h6e;
		memory[16'h1013] <= 8'h27;
		memory[16'h1014] <= 8'hae;
		memory[16'h1015] <= 8'h42;
		memory[16'h1016] <= 8'hc4;
		memory[16'h1017] <= 8'hd8;
		memory[16'h1018] <= 8'h29;
		memory[16'h1019] <= 8'h85;
		memory[16'h101a] <= 8'h75;
		memory[16'h101b] <= 8'h68;
		memory[16'h101c] <= 8'h13;
		memory[16'h101d] <= 8'h41;
		memory[16'h101e] <= 8'h5d;
		memory[16'h101f] <= 8'hc5;
		memory[16'h1020] <= 8'h15;
		memory[16'h1021] <= 8'hb5;
		memory[16'h1022] <= 8'h1e;
		memory[16'h1023] <= 8'hef;
		memory[16'h1024] <= 8'h8e;
		memory[16'h1025] <= 8'hd2;
		memory[16'h1026] <= 8'h4a;
		memory[16'h1027] <= 8'ha6;
		memory[16'h1028] <= 8'h30;
		memory[16'h1029] <= 8'he9;
		memory[16'h102a] <= 8'he6;
		memory[16'h102b] <= 8'he9;
		memory[16'h102c] <= 8'h4d;
		memory[16'h102d] <= 8'had;
		memory[16'h102e] <= 8'h3b;
		memory[16'h102f] <= 8'h31;
		memory[16'h1030] <= 8'h64;
		memory[16'h1031] <= 8'ha9;
		memory[16'h1032] <= 8'h59;
		memory[16'h1033] <= 8'h13;
		memory[16'h1034] <= 8'hec;
		memory[16'h1035] <= 8'h1d;
		memory[16'h1036] <= 8'heb;
		memory[16'h1037] <= 8'h15;
		memory[16'h1038] <= 8'ha3;
		memory[16'h1039] <= 8'h60;
		memory[16'h103a] <= 8'h7d;
		memory[16'h103b] <= 8'hb6;
		memory[16'h103c] <= 8'ha1;
		memory[16'h103d] <= 8'hdb;
		memory[16'h103e] <= 8'h7b;
		memory[16'h103f] <= 8'hb7;
		memory[16'h1040] <= 8'h90;
		memory[16'h1041] <= 8'h9a;
		memory[16'h1042] <= 8'ha6;
		memory[16'h1043] <= 8'h1e;
		memory[16'h1044] <= 8'h6c;
		memory[16'h1045] <= 8'hf0;
		memory[16'h1046] <= 8'hc5;
		memory[16'h1047] <= 8'h9c;
		memory[16'h1048] <= 8'hda;
		memory[16'h1049] <= 8'hab;
		memory[16'h104a] <= 8'h85;
		memory[16'h104b] <= 8'h27;
		memory[16'h104c] <= 8'h59;
		memory[16'h104d] <= 8'hc0;
		memory[16'h104e] <= 8'h59;
		memory[16'h104f] <= 8'hbd;
		memory[16'h1050] <= 8'h6a;
		memory[16'h1051] <= 8'hb2;
		memory[16'h1052] <= 8'hd0;
		memory[16'h1053] <= 8'h56;
		memory[16'h1054] <= 8'hcf;
		memory[16'h1055] <= 8'hbb;
		memory[16'h1056] <= 8'h6b;
		memory[16'h1057] <= 8'h72;
		memory[16'h1058] <= 8'h1c;
		memory[16'h1059] <= 8'he8;
		memory[16'h105a] <= 8'h29;
		memory[16'h105b] <= 8'hbd;
		memory[16'h105c] <= 8'hc3;
		memory[16'h105d] <= 8'ha4;
		memory[16'h105e] <= 8'h74;
		memory[16'h105f] <= 8'h54;
		memory[16'h1060] <= 8'h3e;
		memory[16'h1061] <= 8'h1b;
		memory[16'h1062] <= 8'h72;
		memory[16'h1063] <= 8'haa;
		memory[16'h1064] <= 8'hb;
		memory[16'h1065] <= 8'h37;
		memory[16'h1066] <= 8'h46;
		memory[16'h1067] <= 8'he5;
		memory[16'h1068] <= 8'he3;
		memory[16'h1069] <= 8'hcc;
		memory[16'h106a] <= 8'hd;
		memory[16'h106b] <= 8'h3c;
		memory[16'h106c] <= 8'h8c;
		memory[16'h106d] <= 8'h66;
		memory[16'h106e] <= 8'hf9;
		memory[16'h106f] <= 8'hf6;
		memory[16'h1070] <= 8'h18;
		memory[16'h1071] <= 8'hca;
		memory[16'h1072] <= 8'h4c;
		memory[16'h1073] <= 8'he7;
		memory[16'h1074] <= 8'h85;
		memory[16'h1075] <= 8'hb7;
		memory[16'h1076] <= 8'h5a;
		memory[16'h1077] <= 8'ha1;
		memory[16'h1078] <= 8'ha0;
		memory[16'h1079] <= 8'h83;
		memory[16'h107a] <= 8'h5f;
		memory[16'h107b] <= 8'h63;
		memory[16'h107c] <= 8'h27;
		memory[16'h107d] <= 8'hd3;
		memory[16'h107e] <= 8'hb7;
		memory[16'h107f] <= 8'h66;
		memory[16'h1080] <= 8'hee;
		memory[16'h1081] <= 8'h2a;
		memory[16'h1082] <= 8'h10;
		memory[16'h1083] <= 8'hfa;
		memory[16'h1084] <= 8'h61;
		memory[16'h1085] <= 8'h57;
		memory[16'h1086] <= 8'hdf;
		memory[16'h1087] <= 8'h44;
		memory[16'h1088] <= 8'h23;
		memory[16'h1089] <= 8'hec;
		memory[16'h108a] <= 8'h80;
		memory[16'h108b] <= 8'haf;
		memory[16'h108c] <= 8'h52;
		memory[16'h108d] <= 8'h7a;
		memory[16'h108e] <= 8'ha6;
		memory[16'h108f] <= 8'h6a;
		memory[16'h1090] <= 8'h44;
		memory[16'h1091] <= 8'hf2;
		memory[16'h1092] <= 8'h52;
		memory[16'h1093] <= 8'hc9;
		memory[16'h1094] <= 8'haa;
		memory[16'h1095] <= 8'hac;
		memory[16'h1096] <= 8'h6b;
		memory[16'h1097] <= 8'h4a;
		memory[16'h1098] <= 8'h2f;
		memory[16'h1099] <= 8'hca;
		memory[16'h109a] <= 8'had;
		memory[16'h109b] <= 8'h56;
		memory[16'h109c] <= 8'h9d;
		memory[16'h109d] <= 8'h65;
		memory[16'h109e] <= 8'hbc;
		memory[16'h109f] <= 8'h8c;
		memory[16'h10a0] <= 8'h8f;
		memory[16'h10a1] <= 8'hcd;
		memory[16'h10a2] <= 8'h86;
		memory[16'h10a3] <= 8'hf0;
		memory[16'h10a4] <= 8'h24;
		memory[16'h10a5] <= 8'h65;
		memory[16'h10a6] <= 8'h35;
		memory[16'h10a7] <= 8'h47;
		memory[16'h10a8] <= 8'h52;
		memory[16'h10a9] <= 8'hb5;
		memory[16'h10aa] <= 8'hf6;
		memory[16'h10ab] <= 8'ha4;
		memory[16'h10ac] <= 8'h2f;
		memory[16'h10ad] <= 8'h9c;
		memory[16'h10ae] <= 8'hf;
		memory[16'h10af] <= 8'h73;
		memory[16'h10b0] <= 8'h8f;
		memory[16'h10b1] <= 8'h61;
		memory[16'h10b2] <= 8'h3d;
		memory[16'h10b3] <= 8'h39;
		memory[16'h10b4] <= 8'hd;
		memory[16'h10b5] <= 8'ha8;
		memory[16'h10b6] <= 8'h83;
		memory[16'h10b7] <= 8'h3c;
		memory[16'h10b8] <= 8'h72;
		memory[16'h10b9] <= 8'h30;
		memory[16'h10ba] <= 8'h92;
		memory[16'h10bb] <= 8'hf;
		memory[16'h10bc] <= 8'h95;
		memory[16'h10bd] <= 8'h4f;
		memory[16'h10be] <= 8'h9b;
		memory[16'h10bf] <= 8'h24;
		memory[16'h10c0] <= 8'h1c;
		memory[16'h10c1] <= 8'h21;
		memory[16'h10c2] <= 8'h15;
		memory[16'h10c3] <= 8'h40;
		memory[16'h10c4] <= 8'h87;
		memory[16'h10c5] <= 8'h4a;
		memory[16'h10c6] <= 8'h87;
		memory[16'h10c7] <= 8'hd9;
		memory[16'h10c8] <= 8'hff;
		memory[16'h10c9] <= 8'h7d;
		memory[16'h10ca] <= 8'h7d;
		memory[16'h10cb] <= 8'h2f;
		memory[16'h10cc] <= 8'h1a;
		memory[16'h10cd] <= 8'h8c;
		memory[16'h10ce] <= 8'ha2;
		memory[16'h10cf] <= 8'ha9;
		memory[16'h10d0] <= 8'hed;
		memory[16'h10d1] <= 8'hdf;
		memory[16'h10d2] <= 8'he2;
		memory[16'h10d3] <= 8'hfa;
		memory[16'h10d4] <= 8'h87;
		memory[16'h10d5] <= 8'h65;
		memory[16'h10d6] <= 8'h36;
		memory[16'h10d7] <= 8'hf9;
		memory[16'h10d8] <= 8'h95;
		memory[16'h10d9] <= 8'hc9;
		memory[16'h10da] <= 8'h9;
		memory[16'h10db] <= 8'h2b;
		memory[16'h10dc] <= 8'h18;
		memory[16'h10dd] <= 8'ha4;
		memory[16'h10de] <= 8'h4f;
		memory[16'h10df] <= 8'h34;
		memory[16'h10e0] <= 8'hc6;
		memory[16'h10e1] <= 8'h64;
		memory[16'h10e2] <= 8'h74;
		memory[16'h10e3] <= 8'h4d;
		memory[16'h10e4] <= 8'hae;
		memory[16'h10e5] <= 8'hfb;
		memory[16'h10e6] <= 8'h26;
		memory[16'h10e7] <= 8'hae;
		memory[16'h10e8] <= 8'h78;
		memory[16'h10e9] <= 8'ha3;
		memory[16'h10ea] <= 8'hdd;
		memory[16'h10eb] <= 8'h92;
		memory[16'h10ec] <= 8'h30;
		memory[16'h10ed] <= 8'h7f;
		memory[16'h10ee] <= 8'h3b;
		memory[16'h10ef] <= 8'h1d;
		memory[16'h10f0] <= 8'h5f;
		memory[16'h10f1] <= 8'h1d;
		memory[16'h10f2] <= 8'h18;
		memory[16'h10f3] <= 8'he6;
		memory[16'h10f4] <= 8'h82;
		memory[16'h10f5] <= 8'h4e;
		memory[16'h10f6] <= 8'he0;
		memory[16'h10f7] <= 8'h18;
		memory[16'h10f8] <= 8'h17;
		memory[16'h10f9] <= 8'he9;
		memory[16'h10fa] <= 8'h43;
		memory[16'h10fb] <= 8'h2f;
		memory[16'h10fc] <= 8'h8d;
		memory[16'h10fd] <= 8'h92;
		memory[16'h10fe] <= 8'h63;
		memory[16'h10ff] <= 8'h53;
		memory[16'h1100] <= 8'hf7;
		memory[16'h1101] <= 8'hd7;
		memory[16'h1102] <= 8'ha0;
		memory[16'h1103] <= 8'ha5;
		memory[16'h1104] <= 8'hd2;
		memory[16'h1105] <= 8'hc6;
		memory[16'h1106] <= 8'h53;
		memory[16'h1107] <= 8'h4b;
		memory[16'h1108] <= 8'h6a;
		memory[16'h1109] <= 8'h30;
		memory[16'h110a] <= 8'hdd;
		memory[16'h110b] <= 8'h9a;
		memory[16'h110c] <= 8'hb0;
		memory[16'h110d] <= 8'h19;
		memory[16'h110e] <= 8'hb7;
		memory[16'h110f] <= 8'hf;
		memory[16'h1110] <= 8'h36;
		memory[16'h1111] <= 8'hcf;
		memory[16'h1112] <= 8'hf5;
		memory[16'h1113] <= 8'hb9;
		memory[16'h1114] <= 8'h1e;
		memory[16'h1115] <= 8'hd5;
		memory[16'h1116] <= 8'hd1;
		memory[16'h1117] <= 8'h35;
		memory[16'h1118] <= 8'hbe;
		memory[16'h1119] <= 8'h14;
		memory[16'h111a] <= 8'h65;
		memory[16'h111b] <= 8'h4c;
		memory[16'h111c] <= 8'ha6;
		memory[16'h111d] <= 8'hc8;
		memory[16'h111e] <= 8'h9f;
		memory[16'h111f] <= 8'h9d;
		memory[16'h1120] <= 8'ha0;
		memory[16'h1121] <= 8'h40;
		memory[16'h1122] <= 8'h43;
		memory[16'h1123] <= 8'h72;
		memory[16'h1124] <= 8'h6;
		memory[16'h1125] <= 8'h96;
		memory[16'h1126] <= 8'hbd;
		memory[16'h1127] <= 8'h70;
		memory[16'h1128] <= 8'hc7;
		memory[16'h1129] <= 8'h9b;
		memory[16'h112a] <= 8'ha;
		memory[16'h112b] <= 8'h77;
		memory[16'h112c] <= 8'hb4;
		memory[16'h112d] <= 8'hc2;
		memory[16'h112e] <= 8'h86;
		memory[16'h112f] <= 8'hea;
		memory[16'h1130] <= 8'h91;
		memory[16'h1131] <= 8'h7b;
		memory[16'h1132] <= 8'ha3;
		memory[16'h1133] <= 8'haf;
		memory[16'h1134] <= 8'h51;
		memory[16'h1135] <= 8'h74;
		memory[16'h1136] <= 8'he5;
		memory[16'h1137] <= 8'hf;
		memory[16'h1138] <= 8'h88;
		memory[16'h1139] <= 8'h4a;
		memory[16'h113a] <= 8'h5b;
		memory[16'h113b] <= 8'h2f;
		memory[16'h113c] <= 8'h12;
		memory[16'h113d] <= 8'hfb;
		memory[16'h113e] <= 8'hcc;
		memory[16'h113f] <= 8'hb2;
		memory[16'h1140] <= 8'h3b;
		memory[16'h1141] <= 8'hf;
		memory[16'h1142] <= 8'h25;
		memory[16'h1143] <= 8'h41;
		memory[16'h1144] <= 8'ha6;
		memory[16'h1145] <= 8'he2;
		memory[16'h1146] <= 8'hb2;
		memory[16'h1147] <= 8'h6d;
		memory[16'h1148] <= 8'h7d;
		memory[16'h1149] <= 8'hbc;
		memory[16'h114a] <= 8'he4;
		memory[16'h114b] <= 8'h31;
		memory[16'h114c] <= 8'h7e;
		memory[16'h114d] <= 8'h6a;
		memory[16'h114e] <= 8'h1c;
		memory[16'h114f] <= 8'h10;
		memory[16'h1150] <= 8'he5;
		memory[16'h1151] <= 8'hbf;
		memory[16'h1152] <= 8'hbf;
		memory[16'h1153] <= 8'h36;
		memory[16'h1154] <= 8'h34;
		memory[16'h1155] <= 8'ha4;
		memory[16'h1156] <= 8'h46;
		memory[16'h1157] <= 8'hbc;
		memory[16'h1158] <= 8'hee;
		memory[16'h1159] <= 8'ha1;
		memory[16'h115a] <= 8'heb;
		memory[16'h115b] <= 8'h1;
		memory[16'h115c] <= 8'h9c;
		memory[16'h115d] <= 8'hb8;
		memory[16'h115e] <= 8'hb3;
		memory[16'h115f] <= 8'hd7;
		memory[16'h1160] <= 8'hc7;
		memory[16'h1161] <= 8'hd8;
		memory[16'h1162] <= 8'h19;
		memory[16'h1163] <= 8'h6d;
		memory[16'h1164] <= 8'hbb;
		memory[16'h1165] <= 8'hcb;
		memory[16'h1166] <= 8'hda;
		memory[16'h1167] <= 8'h38;
		memory[16'h1168] <= 8'h87;
		memory[16'h1169] <= 8'hbe;
		memory[16'h116a] <= 8'h6a;
		memory[16'h116b] <= 8'h6;
		memory[16'h116c] <= 8'h28;
		memory[16'h116d] <= 8'h86;
		memory[16'h116e] <= 8'h16;
		memory[16'h116f] <= 8'he;
		memory[16'h1170] <= 8'h45;
		memory[16'h1171] <= 8'hd5;
		memory[16'h1172] <= 8'h44;
		memory[16'h1173] <= 8'h79;
		memory[16'h1174] <= 8'h7a;
		memory[16'h1175] <= 8'h8a;
		memory[16'h1176] <= 8'h36;
		memory[16'h1177] <= 8'h68;
		memory[16'h1178] <= 8'h2c;
		memory[16'h1179] <= 8'h21;
		memory[16'h117a] <= 8'h69;
		memory[16'h117b] <= 8'hc8;
		memory[16'h117c] <= 8'hd9;
		memory[16'h117d] <= 8'h1d;
		memory[16'h117e] <= 8'ha0;
		memory[16'h117f] <= 8'ha1;
		memory[16'h1180] <= 8'hf5;
		memory[16'h1181] <= 8'hb9;
		memory[16'h1182] <= 8'he;
		memory[16'h1183] <= 8'hb0;
		memory[16'h1184] <= 8'h84;
		memory[16'h1185] <= 8'he9;
		memory[16'h1186] <= 8'he9;
		memory[16'h1187] <= 8'hb;
		memory[16'h1188] <= 8'ha7;
		memory[16'h1189] <= 8'h53;
		memory[16'h118a] <= 8'h11;
		memory[16'h118b] <= 8'hd0;
		memory[16'h118c] <= 8'hd9;
		memory[16'h118d] <= 8'h27;
		memory[16'h118e] <= 8'hde;
		memory[16'h118f] <= 8'h1e;
		memory[16'h1190] <= 8'hfd;
		memory[16'h1191] <= 8'h22;
		memory[16'h1192] <= 8'h98;
		memory[16'h1193] <= 8'h77;
		memory[16'h1194] <= 8'had;
		memory[16'h1195] <= 8'hce;
		memory[16'h1196] <= 8'hdf;
		memory[16'h1197] <= 8'hd9;
		memory[16'h1198] <= 8'hef;
		memory[16'h1199] <= 8'h49;
		memory[16'h119a] <= 8'ha1;
		memory[16'h119b] <= 8'hc9;
		memory[16'h119c] <= 8'h66;
		memory[16'h119d] <= 8'h41;
		memory[16'h119e] <= 8'h6a;
		memory[16'h119f] <= 8'h5b;
		memory[16'h11a0] <= 8'hfa;
		memory[16'h11a1] <= 8'h78;
		memory[16'h11a2] <= 8'hc;
		memory[16'h11a3] <= 8'h7e;
		memory[16'h11a4] <= 8'h61;
		memory[16'h11a5] <= 8'hf5;
		memory[16'h11a6] <= 8'h8a;
		memory[16'h11a7] <= 8'h9;
		memory[16'h11a8] <= 8'h48;
		memory[16'h11a9] <= 8'h9b;
		memory[16'h11aa] <= 8'hd9;
		memory[16'h11ab] <= 8'h21;
		memory[16'h11ac] <= 8'hc3;
		memory[16'h11ad] <= 8'hb7;
		memory[16'h11ae] <= 8'h3f;
		memory[16'h11af] <= 8'hc0;
		memory[16'h11b0] <= 8'hd9;
		memory[16'h11b1] <= 8'hd7;
		memory[16'h11b2] <= 8'h37;
		memory[16'h11b3] <= 8'h86;
		memory[16'h11b4] <= 8'ha5;
		memory[16'h11b5] <= 8'h16;
		memory[16'h11b6] <= 8'h5f;
		memory[16'h11b7] <= 8'h95;
		memory[16'h11b8] <= 8'h5f;
		memory[16'h11b9] <= 8'h1;
		memory[16'h11ba] <= 8'h5e;
		memory[16'h11bb] <= 8'hc5;
		memory[16'h11bc] <= 8'h42;
		memory[16'h11bd] <= 8'hc8;
		memory[16'h11be] <= 8'h21;
		memory[16'h11bf] <= 8'h3d;
		memory[16'h11c0] <= 8'h40;
		memory[16'h11c1] <= 8'h2d;
		memory[16'h11c2] <= 8'hbb;
		memory[16'h11c3] <= 8'ha2;
		memory[16'h11c4] <= 8'h22;
		memory[16'h11c5] <= 8'h45;
		memory[16'h11c6] <= 8'hab;
		memory[16'h11c7] <= 8'h6a;
		memory[16'h11c8] <= 8'he1;
		memory[16'h11c9] <= 8'h84;
		memory[16'h11ca] <= 8'h8b;
		memory[16'h11cb] <= 8'ha4;
		memory[16'h11cc] <= 8'h3b;
		memory[16'h11cd] <= 8'hca;
		memory[16'h11ce] <= 8'h64;
		memory[16'h11cf] <= 8'h14;
		memory[16'h11d0] <= 8'ha2;
		memory[16'h11d1] <= 8'h9b;
		memory[16'h11d2] <= 8'h9b;
		memory[16'h11d3] <= 8'h47;
		memory[16'h11d4] <= 8'hb1;
		memory[16'h11d5] <= 8'hfa;
		memory[16'h11d6] <= 8'hdc;
		memory[16'h11d7] <= 8'h11;
		memory[16'h11d8] <= 8'hfb;
		memory[16'h11d9] <= 8'h3a;
		memory[16'h11da] <= 8'hd6;
		memory[16'h11db] <= 8'h3e;
		memory[16'h11dc] <= 8'h2;
		memory[16'h11dd] <= 8'hf7;
		memory[16'h11de] <= 8'h7b;
		memory[16'h11df] <= 8'h43;
		memory[16'h11e0] <= 8'h24;
		memory[16'h11e1] <= 8'h36;
		memory[16'h11e2] <= 8'he5;
		memory[16'h11e3] <= 8'h46;
		memory[16'h11e4] <= 8'h7c;
		memory[16'h11e5] <= 8'h90;
		memory[16'h11e6] <= 8'hb0;
		memory[16'h11e7] <= 8'h5d;
		memory[16'h11e8] <= 8'h14;
		memory[16'h11e9] <= 8'h3b;
		memory[16'h11ea] <= 8'h1;
		memory[16'h11eb] <= 8'h4f;
		memory[16'h11ec] <= 8'h6;
		memory[16'h11ed] <= 8'h65;
		memory[16'h11ee] <= 8'h63;
		memory[16'h11ef] <= 8'ha8;
		memory[16'h11f0] <= 8'h0;
		memory[16'h11f1] <= 8'hfe;
		memory[16'h11f2] <= 8'hef;
		memory[16'h11f3] <= 8'hb1;
		memory[16'h11f4] <= 8'hf9;
		memory[16'h11f5] <= 8'hcc;
		memory[16'h11f6] <= 8'hc2;
		memory[16'h11f7] <= 8'hf4;
		memory[16'h11f8] <= 8'h6;
		memory[16'h11f9] <= 8'h99;
		memory[16'h11fa] <= 8'h32;
		memory[16'h11fb] <= 8'h9;
		memory[16'h11fc] <= 8'h90;
		memory[16'h11fd] <= 8'had;
		memory[16'h11fe] <= 8'h4c;
		memory[16'h11ff] <= 8'hb5;
		memory[16'h1200] <= 8'he4;
		memory[16'h1201] <= 8'h31;
		memory[16'h1202] <= 8'hfb;
		memory[16'h1203] <= 8'h60;
		memory[16'h1204] <= 8'hc1;
		memory[16'h1205] <= 8'hac;
		memory[16'h1206] <= 8'hbd;
		memory[16'h1207] <= 8'hd5;
		memory[16'h1208] <= 8'he7;
		memory[16'h1209] <= 8'hbe;
		memory[16'h120a] <= 8'h24;
		memory[16'h120b] <= 8'hed;
		memory[16'h120c] <= 8'h23;
		memory[16'h120d] <= 8'h87;
		memory[16'h120e] <= 8'h95;
		memory[16'h120f] <= 8'h23;
		memory[16'h1210] <= 8'h86;
		memory[16'h1211] <= 8'h85;
		memory[16'h1212] <= 8'hd4;
		memory[16'h1213] <= 8'h7f;
		memory[16'h1214] <= 8'h51;
		memory[16'h1215] <= 8'h97;
		memory[16'h1216] <= 8'h73;
		memory[16'h1217] <= 8'h57;
		memory[16'h1218] <= 8'h30;
		memory[16'h1219] <= 8'ha6;
		memory[16'h121a] <= 8'h60;
		memory[16'h121b] <= 8'hc0;
		memory[16'h121c] <= 8'h53;
		memory[16'h121d] <= 8'hac;
		memory[16'h121e] <= 8'h75;
		memory[16'h121f] <= 8'h37;
		memory[16'h1220] <= 8'hdd;
		memory[16'h1221] <= 8'h71;
		memory[16'h1222] <= 8'h97;
		memory[16'h1223] <= 8'h9e;
		memory[16'h1224] <= 8'h1d;
		memory[16'h1225] <= 8'h54;
		memory[16'h1226] <= 8'h73;
		memory[16'h1227] <= 8'h4;
		memory[16'h1228] <= 8'h12;
		memory[16'h1229] <= 8'h97;
		memory[16'h122a] <= 8'hf2;
		memory[16'h122b] <= 8'h35;
		memory[16'h122c] <= 8'h1f;
		memory[16'h122d] <= 8'h87;
		memory[16'h122e] <= 8'h58;
		memory[16'h122f] <= 8'ha5;
		memory[16'h1230] <= 8'hc;
		memory[16'h1231] <= 8'h2d;
		memory[16'h1232] <= 8'h24;
		memory[16'h1233] <= 8'h5d;
		memory[16'h1234] <= 8'hc4;
		memory[16'h1235] <= 8'h97;
		memory[16'h1236] <= 8'hb5;
		memory[16'h1237] <= 8'hf4;
		memory[16'h1238] <= 8'h3d;
		memory[16'h1239] <= 8'h15;
		memory[16'h123a] <= 8'hb4;
		memory[16'h123b] <= 8'h91;
		memory[16'h123c] <= 8'hc2;
		memory[16'h123d] <= 8'h2a;
		memory[16'h123e] <= 8'hc8;
		memory[16'h123f] <= 8'h9f;
		memory[16'h1240] <= 8'h9b;
		memory[16'h1241] <= 8'h60;
		memory[16'h1242] <= 8'h3e;
		memory[16'h1243] <= 8'hb8;
		memory[16'h1244] <= 8'hb4;
		memory[16'h1245] <= 8'hb1;
		memory[16'h1246] <= 8'hbc;
		memory[16'h1247] <= 8'hc7;
		memory[16'h1248] <= 8'h49;
		memory[16'h1249] <= 8'hae;
		memory[16'h124a] <= 8'hfc;
		memory[16'h124b] <= 8'h68;
		memory[16'h124c] <= 8'h36;
		memory[16'h124d] <= 8'h55;
		memory[16'h124e] <= 8'hd;
		memory[16'h124f] <= 8'h42;
		memory[16'h1250] <= 8'h82;
		memory[16'h1251] <= 8'h31;
		memory[16'h1252] <= 8'ha0;
		memory[16'h1253] <= 8'h46;
		memory[16'h1254] <= 8'hc8;
		memory[16'h1255] <= 8'h55;
		memory[16'h1256] <= 8'h3a;
		memory[16'h1257] <= 8'h6;
		memory[16'h1258] <= 8'h6a;
		memory[16'h1259] <= 8'hee;
		memory[16'h125a] <= 8'h97;
		memory[16'h125b] <= 8'h2c;
		memory[16'h125c] <= 8'h18;
		memory[16'h125d] <= 8'h5f;
		memory[16'h125e] <= 8'hcc;
		memory[16'h125f] <= 8'hb3;
		memory[16'h1260] <= 8'hbf;
		memory[16'h1261] <= 8'ha;
		memory[16'h1262] <= 8'h6b;
		memory[16'h1263] <= 8'h74;
		memory[16'h1264] <= 8'hbb;
		memory[16'h1265] <= 8'h28;
		memory[16'h1266] <= 8'h3b;
		memory[16'h1267] <= 8'h4;
		memory[16'h1268] <= 8'hd6;
		memory[16'h1269] <= 8'h37;
		memory[16'h126a] <= 8'h6c;
		memory[16'h126b] <= 8'hc;
		memory[16'h126c] <= 8'h8c;
		memory[16'h126d] <= 8'h79;
		memory[16'h126e] <= 8'h4f;
		memory[16'h126f] <= 8'he;
		memory[16'h1270] <= 8'haa;
		memory[16'h1271] <= 8'hef;
		memory[16'h1272] <= 8'h54;
		memory[16'h1273] <= 8'h73;
		memory[16'h1274] <= 8'h44;
		memory[16'h1275] <= 8'h8e;
		memory[16'h1276] <= 8'h79;
		memory[16'h1277] <= 8'hae;
		memory[16'h1278] <= 8'h7d;
		memory[16'h1279] <= 8'h10;
		memory[16'h127a] <= 8'hdb;
		memory[16'h127b] <= 8'h95;
		memory[16'h127c] <= 8'h6f;
		memory[16'h127d] <= 8'ha7;
		memory[16'h127e] <= 8'h49;
		memory[16'h127f] <= 8'h2f;
		memory[16'h1280] <= 8'hb1;
		memory[16'h1281] <= 8'hb4;
		memory[16'h1282] <= 8'ha3;
		memory[16'h1283] <= 8'h6c;
		memory[16'h1284] <= 8'hdc;
		memory[16'h1285] <= 8'hde;
		memory[16'h1286] <= 8'h71;
		memory[16'h1287] <= 8'hb3;
		memory[16'h1288] <= 8'h15;
		memory[16'h1289] <= 8'hdd;
		memory[16'h128a] <= 8'hbf;
		memory[16'h128b] <= 8'ha2;
		memory[16'h128c] <= 8'h57;
		memory[16'h128d] <= 8'he;
		memory[16'h128e] <= 8'hb0;
		memory[16'h128f] <= 8'h1;
		memory[16'h1290] <= 8'hfd;
		memory[16'h1291] <= 8'h5;
		memory[16'h1292] <= 8'h74;
		memory[16'h1293] <= 8'h41;
		memory[16'h1294] <= 8'h93;
		memory[16'h1295] <= 8'hed;
		memory[16'h1296] <= 8'hf0;
		memory[16'h1297] <= 8'h10;
		memory[16'h1298] <= 8'hfd;
		memory[16'h1299] <= 8'hcb;
		memory[16'h129a] <= 8'ha6;
		memory[16'h129b] <= 8'h6d;
		memory[16'h129c] <= 8'h72;
		memory[16'h129d] <= 8'hef;
		memory[16'h129e] <= 8'h9c;
		memory[16'h129f] <= 8'h23;
		memory[16'h12a0] <= 8'ha3;
		memory[16'h12a1] <= 8'h3f;
		memory[16'h12a2] <= 8'h8f;
		memory[16'h12a3] <= 8'h80;
		memory[16'h12a4] <= 8'h1d;
		memory[16'h12a5] <= 8'h0;
		memory[16'h12a6] <= 8'h33;
		memory[16'h12a7] <= 8'h32;
		memory[16'h12a8] <= 8'hde;
		memory[16'h12a9] <= 8'hf2;
		memory[16'h12aa] <= 8'hd4;
		memory[16'h12ab] <= 8'h35;
		memory[16'h12ac] <= 8'h1;
		memory[16'h12ad] <= 8'h85;
		memory[16'h12ae] <= 8'h36;
		memory[16'h12af] <= 8'hfe;
		memory[16'h12b0] <= 8'h8a;
		memory[16'h12b1] <= 8'hab;
		memory[16'h12b2] <= 8'h40;
		memory[16'h12b3] <= 8'h1d;
		memory[16'h12b4] <= 8'h98;
		memory[16'h12b5] <= 8'h30;
		memory[16'h12b6] <= 8'h2e;
		memory[16'h12b7] <= 8'h96;
		memory[16'h12b8] <= 8'hfb;
		memory[16'h12b9] <= 8'hd4;
		memory[16'h12ba] <= 8'h3;
		memory[16'h12bb] <= 8'h6d;
		memory[16'h12bc] <= 8'hc3;
		memory[16'h12bd] <= 8'h9f;
		memory[16'h12be] <= 8'h90;
		memory[16'h12bf] <= 8'h66;
		memory[16'h12c0] <= 8'hde;
		memory[16'h12c1] <= 8'h1f;
		memory[16'h12c2] <= 8'he6;
		memory[16'h12c3] <= 8'hfb;
		memory[16'h12c4] <= 8'h20;
		memory[16'h12c5] <= 8'h19;
		memory[16'h12c6] <= 8'h2d;
		memory[16'h12c7] <= 8'hfe;
		memory[16'h12c8] <= 8'hc;
		memory[16'h12c9] <= 8'h2;
		memory[16'h12ca] <= 8'h33;
		memory[16'h12cb] <= 8'hd;
		memory[16'h12cc] <= 8'h87;
		memory[16'h12cd] <= 8'h69;
		memory[16'h12ce] <= 8'hb;
		memory[16'h12cf] <= 8'h11;
		memory[16'h12d0] <= 8'h14;
		memory[16'h12d1] <= 8'h4b;
		memory[16'h12d2] <= 8'h2e;
		memory[16'h12d3] <= 8'had;
		memory[16'h12d4] <= 8'h7b;
		memory[16'h12d5] <= 8'h5c;
		memory[16'h12d6] <= 8'h43;
		memory[16'h12d7] <= 8'h76;
		memory[16'h12d8] <= 8'h30;
		memory[16'h12d9] <= 8'h46;
		memory[16'h12da] <= 8'he3;
		memory[16'h12db] <= 8'hf3;
		memory[16'h12dc] <= 8'he5;
		memory[16'h12dd] <= 8'h73;
		memory[16'h12de] <= 8'h5a;
		memory[16'h12df] <= 8'hc3;
		memory[16'h12e0] <= 8'h93;
		memory[16'h12e1] <= 8'h40;
		memory[16'h12e2] <= 8'hbe;
		memory[16'h12e3] <= 8'hb3;
		memory[16'h12e4] <= 8'h5a;
		memory[16'h12e5] <= 8'heb;
		memory[16'h12e6] <= 8'hb1;
		memory[16'h12e7] <= 8'h66;
		memory[16'h12e8] <= 8'hed;
		memory[16'h12e9] <= 8'he4;
		memory[16'h12ea] <= 8'h73;
		memory[16'h12eb] <= 8'h74;
		memory[16'h12ec] <= 8'h4d;
		memory[16'h12ed] <= 8'h7e;
		memory[16'h12ee] <= 8'h85;
		memory[16'h12ef] <= 8'h62;
		memory[16'h12f0] <= 8'hca;
		memory[16'h12f1] <= 8'hb4;
		memory[16'h12f2] <= 8'hf;
		memory[16'h12f3] <= 8'h45;
		memory[16'h12f4] <= 8'h10;
		memory[16'h12f5] <= 8'h52;
		memory[16'h12f6] <= 8'hbc;
		memory[16'h12f7] <= 8'h41;
		memory[16'h12f8] <= 8'h98;
		memory[16'h12f9] <= 8'h9f;
		memory[16'h12fa] <= 8'h34;
		memory[16'h12fb] <= 8'h7d;
		memory[16'h12fc] <= 8'h13;
		memory[16'h12fd] <= 8'h8e;
		memory[16'h12fe] <= 8'h40;
		memory[16'h12ff] <= 8'ha6;
		memory[16'h1300] <= 8'hcf;
		memory[16'h1301] <= 8'hfe;
		memory[16'h1302] <= 8'h59;
		memory[16'h1303] <= 8'h29;
		memory[16'h1304] <= 8'he9;
		memory[16'h1305] <= 8'ha;
		memory[16'h1306] <= 8'h8f;
		memory[16'h1307] <= 8'hd7;
		memory[16'h1308] <= 8'hee;
		memory[16'h1309] <= 8'h2;
		memory[16'h130a] <= 8'h4b;
		memory[16'h130b] <= 8'h3b;
		memory[16'h130c] <= 8'h80;
		memory[16'h130d] <= 8'hd1;
		memory[16'h130e] <= 8'h9d;
		memory[16'h130f] <= 8'h4a;
		memory[16'h1310] <= 8'h85;
		memory[16'h1311] <= 8'hac;
		memory[16'h1312] <= 8'h90;
		memory[16'h1313] <= 8'h95;
		memory[16'h1314] <= 8'hfe;
		memory[16'h1315] <= 8'h4c;
		memory[16'h1316] <= 8'hd6;
		memory[16'h1317] <= 8'h96;
		memory[16'h1318] <= 8'heb;
		memory[16'h1319] <= 8'hb;
		memory[16'h131a] <= 8'h13;
		memory[16'h131b] <= 8'hfe;
		memory[16'h131c] <= 8'h99;
		memory[16'h131d] <= 8'h53;
		memory[16'h131e] <= 8'ha4;
		memory[16'h131f] <= 8'h68;
		memory[16'h1320] <= 8'h51;
		memory[16'h1321] <= 8'hfd;
		memory[16'h1322] <= 8'h91;
		memory[16'h1323] <= 8'h3b;
		memory[16'h1324] <= 8'h7;
		memory[16'h1325] <= 8'h20;
		memory[16'h1326] <= 8'h12;
		memory[16'h1327] <= 8'hf5;
		memory[16'h1328] <= 8'h22;
		memory[16'h1329] <= 8'h5d;
		memory[16'h132a] <= 8'h31;
		memory[16'h132b] <= 8'ha3;
		memory[16'h132c] <= 8'h2e;
		memory[16'h132d] <= 8'hce;
		memory[16'h132e] <= 8'hed;
		memory[16'h132f] <= 8'hb3;
		memory[16'h1330] <= 8'h7b;
		memory[16'h1331] <= 8'h7d;
		memory[16'h1332] <= 8'h49;
		memory[16'h1333] <= 8'h79;
		memory[16'h1334] <= 8'hc9;
		memory[16'h1335] <= 8'h1f;
		memory[16'h1336] <= 8'h10;
		memory[16'h1337] <= 8'hb5;
		memory[16'h1338] <= 8'h2a;
		memory[16'h1339] <= 8'h23;
		memory[16'h133a] <= 8'hb3;
		memory[16'h133b] <= 8'hc4;
		memory[16'h133c] <= 8'h77;
		memory[16'h133d] <= 8'h58;
		memory[16'h133e] <= 8'h2c;
		memory[16'h133f] <= 8'hc8;
		memory[16'h1340] <= 8'h55;
		memory[16'h1341] <= 8'hbe;
		memory[16'h1342] <= 8'h3;
		memory[16'h1343] <= 8'h5d;
		memory[16'h1344] <= 8'hde;
		memory[16'h1345] <= 8'h15;
		memory[16'h1346] <= 8'h52;
		memory[16'h1347] <= 8'h1;
		memory[16'h1348] <= 8'h73;
		memory[16'h1349] <= 8'h83;
		memory[16'h134a] <= 8'ha4;
		memory[16'h134b] <= 8'ha1;
		memory[16'h134c] <= 8'h52;
		memory[16'h134d] <= 8'h91;
		memory[16'h134e] <= 8'h55;
		memory[16'h134f] <= 8'hcd;
		memory[16'h1350] <= 8'hf;
		memory[16'h1351] <= 8'h9e;
		memory[16'h1352] <= 8'h46;
		memory[16'h1353] <= 8'hd8;
		memory[16'h1354] <= 8'hbd;
		memory[16'h1355] <= 8'h56;
		memory[16'h1356] <= 8'h8d;
		memory[16'h1357] <= 8'he8;
		memory[16'h1358] <= 8'h7a;
		memory[16'h1359] <= 8'h41;
		memory[16'h135a] <= 8'hac;
		memory[16'h135b] <= 8'hf1;
		memory[16'h135c] <= 8'h99;
		memory[16'h135d] <= 8'hd8;
		memory[16'h135e] <= 8'hb9;
		memory[16'h135f] <= 8'hee;
		memory[16'h1360] <= 8'h96;
		memory[16'h1361] <= 8'hbd;
		memory[16'h1362] <= 8'h4b;
		memory[16'h1363] <= 8'h75;
		memory[16'h1364] <= 8'hd2;
		memory[16'h1365] <= 8'h9e;
		memory[16'h1366] <= 8'h76;
		memory[16'h1367] <= 8'h45;
		memory[16'h1368] <= 8'h21;
		memory[16'h1369] <= 8'h1a;
		memory[16'h136a] <= 8'he7;
		memory[16'h136b] <= 8'h73;
		memory[16'h136c] <= 8'hab;
		memory[16'h136d] <= 8'h3c;
		memory[16'h136e] <= 8'h40;
		memory[16'h136f] <= 8'hba;
		memory[16'h1370] <= 8'hda;
		memory[16'h1371] <= 8'h87;
		memory[16'h1372] <= 8'h93;
		memory[16'h1373] <= 8'h97;
		memory[16'h1374] <= 8'hdd;
		memory[16'h1375] <= 8'h20;
		memory[16'h1376] <= 8'h7f;
		memory[16'h1377] <= 8'h57;
		memory[16'h1378] <= 8'h61;
		memory[16'h1379] <= 8'h2b;
		memory[16'h137a] <= 8'h48;
		memory[16'h137b] <= 8'hfa;
		memory[16'h137c] <= 8'h4;
		memory[16'h137d] <= 8'h2;
		memory[16'h137e] <= 8'he9;
		memory[16'h137f] <= 8'h9a;
		memory[16'h1380] <= 8'hbf;
		memory[16'h1381] <= 8'h34;
		memory[16'h1382] <= 8'hf;
		memory[16'h1383] <= 8'h91;
		memory[16'h1384] <= 8'hd2;
		memory[16'h1385] <= 8'h85;
		memory[16'h1386] <= 8'hd7;
		memory[16'h1387] <= 8'hf4;
		memory[16'h1388] <= 8'h9f;
		memory[16'h1389] <= 8'hbe;
		memory[16'h138a] <= 8'h67;
		memory[16'h138b] <= 8'h4b;
		memory[16'h138c] <= 8'hfa;
		memory[16'h138d] <= 8'ha8;
		memory[16'h138e] <= 8'h5;
		memory[16'h138f] <= 8'hd4;
		memory[16'h1390] <= 8'h2f;
		memory[16'h1391] <= 8'h98;
		memory[16'h1392] <= 8'h6b;
		memory[16'h1393] <= 8'hc;
		memory[16'h1394] <= 8'hb9;
		memory[16'h1395] <= 8'heb;
		memory[16'h1396] <= 8'h64;
		memory[16'h1397] <= 8'h1a;
		memory[16'h1398] <= 8'h16;
		memory[16'h1399] <= 8'hac;
		memory[16'h139a] <= 8'h15;
		memory[16'h139b] <= 8'h1a;
		memory[16'h139c] <= 8'hae;
		memory[16'h139d] <= 8'hfe;
		memory[16'h139e] <= 8'hb5;
		memory[16'h139f] <= 8'h6d;
		memory[16'h13a0] <= 8'h32;
		memory[16'h13a1] <= 8'hc4;
		memory[16'h13a2] <= 8'hff;
		memory[16'h13a3] <= 8'h5;
		memory[16'h13a4] <= 8'h4a;
		memory[16'h13a5] <= 8'hd6;
		memory[16'h13a6] <= 8'hf9;
		memory[16'h13a7] <= 8'he9;
		memory[16'h13a8] <= 8'h94;
		memory[16'h13a9] <= 8'h60;
		memory[16'h13aa] <= 8'h34;
		memory[16'h13ab] <= 8'h8e;
		memory[16'h13ac] <= 8'h8;
		memory[16'h13ad] <= 8'h3a;
		memory[16'h13ae] <= 8'h62;
		memory[16'h13af] <= 8'h37;
		memory[16'h13b0] <= 8'hd2;
		memory[16'h13b1] <= 8'hcd;
		memory[16'h13b2] <= 8'h44;
		memory[16'h13b3] <= 8'h8b;
		memory[16'h13b4] <= 8'hb8;
		memory[16'h13b5] <= 8'ha8;
		memory[16'h13b6] <= 8'ha6;
		memory[16'h13b7] <= 8'hcf;
		memory[16'h13b8] <= 8'h54;
		memory[16'h13b9] <= 8'hbb;
		memory[16'h13ba] <= 8'he9;
		memory[16'h13bb] <= 8'h3;
		memory[16'h13bc] <= 8'hb9;
		memory[16'h13bd] <= 8'h9e;
		memory[16'h13be] <= 8'h70;
		memory[16'h13bf] <= 8'heb;
		memory[16'h13c0] <= 8'h63;
		memory[16'h13c1] <= 8'h6f;
		memory[16'h13c2] <= 8'hf0;
		memory[16'h13c3] <= 8'had;
		memory[16'h13c4] <= 8'h45;
		memory[16'h13c5] <= 8'he9;
		memory[16'h13c6] <= 8'h96;
		memory[16'h13c7] <= 8'hd9;
		memory[16'h13c8] <= 8'h4a;
		memory[16'h13c9] <= 8'hcb;
		memory[16'h13ca] <= 8'h67;
		memory[16'h13cb] <= 8'h52;
		memory[16'h13cc] <= 8'h5;
		memory[16'h13cd] <= 8'hc9;
		memory[16'h13ce] <= 8'h8a;
		memory[16'h13cf] <= 8'hd7;
		memory[16'h13d0] <= 8'h97;
		memory[16'h13d1] <= 8'hce;
		memory[16'h13d2] <= 8'h63;
		memory[16'h13d3] <= 8'h4f;
		memory[16'h13d4] <= 8'h76;
		memory[16'h13d5] <= 8'h9;
		memory[16'h13d6] <= 8'h1e;
		memory[16'h13d7] <= 8'hca;
		memory[16'h13d8] <= 8'hc4;
		memory[16'h13d9] <= 8'h8;
		memory[16'h13da] <= 8'hcd;
		memory[16'h13db] <= 8'h7d;
		memory[16'h13dc] <= 8'ha6;
		memory[16'h13dd] <= 8'h3e;
		memory[16'h13de] <= 8'h68;
		memory[16'h13df] <= 8'h9;
		memory[16'h13e0] <= 8'had;
		memory[16'h13e1] <= 8'h59;
		memory[16'h13e2] <= 8'hb6;
		memory[16'h13e3] <= 8'hf3;
		memory[16'h13e4] <= 8'h42;
		memory[16'h13e5] <= 8'h4d;
		memory[16'h13e6] <= 8'hcc;
		memory[16'h13e7] <= 8'h8c;
		memory[16'h13e8] <= 8'h18;
		memory[16'h13e9] <= 8'h34;
		memory[16'h13ea] <= 8'hdf;
		memory[16'h13eb] <= 8'h1d;
		memory[16'h13ec] <= 8'hfd;
		memory[16'h13ed] <= 8'h69;
		memory[16'h13ee] <= 8'hf4;
		memory[16'h13ef] <= 8'h94;
		memory[16'h13f0] <= 8'h37;
		memory[16'h13f1] <= 8'h57;
		memory[16'h13f2] <= 8'he4;
		memory[16'h13f3] <= 8'had;
		memory[16'h13f4] <= 8'h60;
		memory[16'h13f5] <= 8'h2;
		memory[16'h13f6] <= 8'h77;
		memory[16'h13f7] <= 8'h24;
		memory[16'h13f8] <= 8'ha;
		memory[16'h13f9] <= 8'h45;
		memory[16'h13fa] <= 8'ha1;
		memory[16'h13fb] <= 8'hb1;
		memory[16'h13fc] <= 8'h83;
		memory[16'h13fd] <= 8'ha;
		memory[16'h13fe] <= 8'hba;
		memory[16'h13ff] <= 8'h30;
		memory[16'h1400] <= 8'h63;
		memory[16'h1401] <= 8'h71;
		memory[16'h1402] <= 8'h23;
		memory[16'h1403] <= 8'ha5;
		memory[16'h1404] <= 8'hbe;
		memory[16'h1405] <= 8'hf0;
		memory[16'h1406] <= 8'h32;
		memory[16'h1407] <= 8'hd6;
		memory[16'h1408] <= 8'h24;
		memory[16'h1409] <= 8'h11;
		memory[16'h140a] <= 8'hf3;
		memory[16'h140b] <= 8'h21;
		memory[16'h140c] <= 8'h7a;
		memory[16'h140d] <= 8'he7;
		memory[16'h140e] <= 8'hb6;
		memory[16'h140f] <= 8'hb1;
		memory[16'h1410] <= 8'h3f;
		memory[16'h1411] <= 8'h9a;
		memory[16'h1412] <= 8'h5e;
		memory[16'h1413] <= 8'h9f;
		memory[16'h1414] <= 8'h9c;
		memory[16'h1415] <= 8'hd5;
		memory[16'h1416] <= 8'hc4;
		memory[16'h1417] <= 8'ha7;
		memory[16'h1418] <= 8'h1a;
		memory[16'h1419] <= 8'h65;
		memory[16'h141a] <= 8'h58;
		memory[16'h141b] <= 8'h9d;
		memory[16'h141c] <= 8'h6f;
		memory[16'h141d] <= 8'h12;
		memory[16'h141e] <= 8'hce;
		memory[16'h141f] <= 8'hd2;
		memory[16'h1420] <= 8'h83;
		memory[16'h1421] <= 8'hf1;
		memory[16'h1422] <= 8'h78;
		memory[16'h1423] <= 8'h41;
		memory[16'h1424] <= 8'he1;
		memory[16'h1425] <= 8'haa;
		memory[16'h1426] <= 8'h17;
		memory[16'h1427] <= 8'h5;
		memory[16'h1428] <= 8'hbb;
		memory[16'h1429] <= 8'ha;
		memory[16'h142a] <= 8'h27;
		memory[16'h142b] <= 8'h35;
		memory[16'h142c] <= 8'hf2;
		memory[16'h142d] <= 8'hdd;
		memory[16'h142e] <= 8'he6;
		memory[16'h142f] <= 8'h31;
		memory[16'h1430] <= 8'h77;
		memory[16'h1431] <= 8'h44;
		memory[16'h1432] <= 8'hd0;
		memory[16'h1433] <= 8'h13;
		memory[16'h1434] <= 8'h19;
		memory[16'h1435] <= 8'h94;
		memory[16'h1436] <= 8'hba;
		memory[16'h1437] <= 8'h34;
		memory[16'h1438] <= 8'hfa;
		memory[16'h1439] <= 8'h12;
		memory[16'h143a] <= 8'hd1;
		memory[16'h143b] <= 8'h69;
		memory[16'h143c] <= 8'h25;
		memory[16'h143d] <= 8'h9f;
		memory[16'h143e] <= 8'h3c;
		memory[16'h143f] <= 8'ha8;
		memory[16'h1440] <= 8'h91;
		memory[16'h1441] <= 8'hb4;
		memory[16'h1442] <= 8'hea;
		memory[16'h1443] <= 8'h72;
		memory[16'h1444] <= 8'h5e;
		memory[16'h1445] <= 8'h1;
		memory[16'h1446] <= 8'h78;
		memory[16'h1447] <= 8'h19;
		memory[16'h1448] <= 8'hc;
		memory[16'h1449] <= 8'h9f;
		memory[16'h144a] <= 8'h4e;
		memory[16'h144b] <= 8'hfe;
		memory[16'h144c] <= 8'h7c;
		memory[16'h144d] <= 8'h34;
		memory[16'h144e] <= 8'h2f;
		memory[16'h144f] <= 8'hf3;
		memory[16'h1450] <= 8'h78;
		memory[16'h1451] <= 8'hff;
		memory[16'h1452] <= 8'h6;
		memory[16'h1453] <= 8'h91;
		memory[16'h1454] <= 8'h94;
		memory[16'h1455] <= 8'hc1;
		memory[16'h1456] <= 8'hc5;
		memory[16'h1457] <= 8'h8e;
		memory[16'h1458] <= 8'hd3;
		memory[16'h1459] <= 8'h97;
		memory[16'h145a] <= 8'hf7;
		memory[16'h145b] <= 8'hf8;
		memory[16'h145c] <= 8'h36;
		memory[16'h145d] <= 8'h33;
		memory[16'h145e] <= 8'ha1;
		memory[16'h145f] <= 8'hc7;
		memory[16'h1460] <= 8'he7;
		memory[16'h1461] <= 8'h8b;
		memory[16'h1462] <= 8'h3a;
		memory[16'h1463] <= 8'h45;
		memory[16'h1464] <= 8'h8c;
		memory[16'h1465] <= 8'hb2;
		memory[16'h1466] <= 8'h5e;
		memory[16'h1467] <= 8'h98;
		memory[16'h1468] <= 8'h51;
		memory[16'h1469] <= 8'hac;
		memory[16'h146a] <= 8'h96;
		memory[16'h146b] <= 8'hcd;
		memory[16'h146c] <= 8'he0;
		memory[16'h146d] <= 8'hc5;
		memory[16'h146e] <= 8'hc0;
		memory[16'h146f] <= 8'h58;
		memory[16'h1470] <= 8'hc5;
		memory[16'h1471] <= 8'hc6;
		memory[16'h1472] <= 8'hea;
		memory[16'h1473] <= 8'h59;
		memory[16'h1474] <= 8'h87;
		memory[16'h1475] <= 8'haf;
		memory[16'h1476] <= 8'he7;
		memory[16'h1477] <= 8'h5b;
		memory[16'h1478] <= 8'h46;
		memory[16'h1479] <= 8'hde;
		memory[16'h147a] <= 8'h53;
		memory[16'h147b] <= 8'h7d;
		memory[16'h147c] <= 8'h12;
		memory[16'h147d] <= 8'hf4;
		memory[16'h147e] <= 8'h44;
		memory[16'h147f] <= 8'hf9;
		memory[16'h1480] <= 8'h7f;
		memory[16'h1481] <= 8'h7e;
		memory[16'h1482] <= 8'h3f;
		memory[16'h1483] <= 8'hc;
		memory[16'h1484] <= 8'h30;
		memory[16'h1485] <= 8'h9d;
		memory[16'h1486] <= 8'ha4;
		memory[16'h1487] <= 8'h81;
		memory[16'h1488] <= 8'h4a;
		memory[16'h1489] <= 8'h3b;
		memory[16'h148a] <= 8'h4e;
		memory[16'h148b] <= 8'h2a;
		memory[16'h148c] <= 8'h0;
		memory[16'h148d] <= 8'he;
		memory[16'h148e] <= 8'h83;
		memory[16'h148f] <= 8'hc5;
		memory[16'h1490] <= 8'hd5;
		memory[16'h1491] <= 8'h6d;
		memory[16'h1492] <= 8'h1e;
		memory[16'h1493] <= 8'h5c;
		memory[16'h1494] <= 8'h1c;
		memory[16'h1495] <= 8'h5;
		memory[16'h1496] <= 8'hb7;
		memory[16'h1497] <= 8'h63;
		memory[16'h1498] <= 8'he4;
		memory[16'h1499] <= 8'hb;
		memory[16'h149a] <= 8'he0;
		memory[16'h149b] <= 8'hf6;
		memory[16'h149c] <= 8'hff;
		memory[16'h149d] <= 8'h24;
		memory[16'h149e] <= 8'hef;
		memory[16'h149f] <= 8'h7f;
		memory[16'h14a0] <= 8'ha3;
		memory[16'h14a1] <= 8'h2e;
		memory[16'h14a2] <= 8'h8b;
		memory[16'h14a3] <= 8'hd3;
		memory[16'h14a4] <= 8'hcc;
		memory[16'h14a5] <= 8'h2f;
		memory[16'h14a6] <= 8'h55;
		memory[16'h14a7] <= 8'h16;
		memory[16'h14a8] <= 8'h6a;
		memory[16'h14a9] <= 8'ha3;
		memory[16'h14aa] <= 8'h40;
		memory[16'h14ab] <= 8'h6b;
		memory[16'h14ac] <= 8'hb2;
		memory[16'h14ad] <= 8'hc3;
		memory[16'h14ae] <= 8'h30;
		memory[16'h14af] <= 8'h87;
		memory[16'h14b0] <= 8'h30;
		memory[16'h14b1] <= 8'h4f;
		memory[16'h14b2] <= 8'he3;
		memory[16'h14b3] <= 8'h4d;
		memory[16'h14b4] <= 8'h54;
		memory[16'h14b5] <= 8'h9b;
		memory[16'h14b6] <= 8'hb0;
		memory[16'h14b7] <= 8'h38;
		memory[16'h14b8] <= 8'ha6;
		memory[16'h14b9] <= 8'h90;
		memory[16'h14ba] <= 8'h2e;
		memory[16'h14bb] <= 8'ha5;
		memory[16'h14bc] <= 8'hb4;
		memory[16'h14bd] <= 8'h1e;
		memory[16'h14be] <= 8'h24;
		memory[16'h14bf] <= 8'h57;
		memory[16'h14c0] <= 8'h4c;
		memory[16'h14c1] <= 8'haf;
		memory[16'h14c2] <= 8'h2b;
		memory[16'h14c3] <= 8'h18;
		memory[16'h14c4] <= 8'hdf;
		memory[16'h14c5] <= 8'h80;
		memory[16'h14c6] <= 8'h2e;
		memory[16'h14c7] <= 8'h49;
		memory[16'h14c8] <= 8'h23;
		memory[16'h14c9] <= 8'h6f;
		memory[16'h14ca] <= 8'hb4;
		memory[16'h14cb] <= 8'hd5;
		memory[16'h14cc] <= 8'h32;
		memory[16'h14cd] <= 8'he5;
		memory[16'h14ce] <= 8'h5c;
		memory[16'h14cf] <= 8'h63;
		memory[16'h14d0] <= 8'h34;
		memory[16'h14d1] <= 8'h40;
		memory[16'h14d2] <= 8'hb0;
		memory[16'h14d3] <= 8'h88;
		memory[16'h14d4] <= 8'hdb;
		memory[16'h14d5] <= 8'h60;
		memory[16'h14d6] <= 8'hc1;
		memory[16'h14d7] <= 8'h81;
		memory[16'h14d8] <= 8'hf0;
		memory[16'h14d9] <= 8'hef;
		memory[16'h14da] <= 8'h26;
		memory[16'h14db] <= 8'ha4;
		memory[16'h14dc] <= 8'hd;
		memory[16'h14dd] <= 8'h4b;
		memory[16'h14de] <= 8'hfc;
		memory[16'h14df] <= 8'h5a;
		memory[16'h14e0] <= 8'hfa;
		memory[16'h14e1] <= 8'h27;
		memory[16'h14e2] <= 8'h72;
		memory[16'h14e3] <= 8'hd9;
		memory[16'h14e4] <= 8'ha7;
		memory[16'h14e5] <= 8'ha1;
		memory[16'h14e6] <= 8'h23;
		memory[16'h14e7] <= 8'hca;
		memory[16'h14e8] <= 8'h10;
		memory[16'h14e9] <= 8'hd7;
		memory[16'h14ea] <= 8'ha0;
		memory[16'h14eb] <= 8'h42;
		memory[16'h14ec] <= 8'hbc;
		memory[16'h14ed] <= 8'hfc;
		memory[16'h14ee] <= 8'ha5;
		memory[16'h14ef] <= 8'hf0;
		memory[16'h14f0] <= 8'h3c;
		memory[16'h14f1] <= 8'h55;
		memory[16'h14f2] <= 8'h79;
		memory[16'h14f3] <= 8'h17;
		memory[16'h14f4] <= 8'hb5;
		memory[16'h14f5] <= 8'h3a;
		memory[16'h14f6] <= 8'h98;
		memory[16'h14f7] <= 8'ha5;
		memory[16'h14f8] <= 8'h29;
		memory[16'h14f9] <= 8'hbf;
		memory[16'h14fa] <= 8'h4a;
		memory[16'h14fb] <= 8'h37;
		memory[16'h14fc] <= 8'ha;
		memory[16'h14fd] <= 8'h46;
		memory[16'h14fe] <= 8'h91;
		memory[16'h14ff] <= 8'h4;
		memory[16'h1500] <= 8'h6d;
		memory[16'h1501] <= 8'h3;
		memory[16'h1502] <= 8'hde;
		memory[16'h1503] <= 8'h14;
		memory[16'h1504] <= 8'ha4;
		memory[16'h1505] <= 8'h1;
		memory[16'h1506] <= 8'hde;
		memory[16'h1507] <= 8'hb4;
		memory[16'h1508] <= 8'hd8;
		memory[16'h1509] <= 8'h7e;
		memory[16'h150a] <= 8'hf7;
		memory[16'h150b] <= 8'h95;
		memory[16'h150c] <= 8'h7b;
		memory[16'h150d] <= 8'h9c;
		memory[16'h150e] <= 8'h85;
		memory[16'h150f] <= 8'hb7;
		memory[16'h1510] <= 8'hf2;
		memory[16'h1511] <= 8'hfe;
		memory[16'h1512] <= 8'hcf;
		memory[16'h1513] <= 8'ha7;
		memory[16'h1514] <= 8'h38;
		memory[16'h1515] <= 8'h67;
		memory[16'h1516] <= 8'h4d;
		memory[16'h1517] <= 8'h62;
		memory[16'h1518] <= 8'h26;
		memory[16'h1519] <= 8'h97;
		memory[16'h151a] <= 8'h99;
		memory[16'h151b] <= 8'h30;
		memory[16'h151c] <= 8'hdd;
		memory[16'h151d] <= 8'h2a;
		memory[16'h151e] <= 8'h35;
		memory[16'h151f] <= 8'h4a;
		memory[16'h1520] <= 8'h2d;
		memory[16'h1521] <= 8'h13;
		memory[16'h1522] <= 8'h5e;
		memory[16'h1523] <= 8'hd2;
		memory[16'h1524] <= 8'h14;
		memory[16'h1525] <= 8'h3c;
		memory[16'h1526] <= 8'h86;
		memory[16'h1527] <= 8'hec;
		memory[16'h1528] <= 8'hbb;
		memory[16'h1529] <= 8'h7d;
		memory[16'h152a] <= 8'h81;
		memory[16'h152b] <= 8'h36;
		memory[16'h152c] <= 8'h1a;
		memory[16'h152d] <= 8'h7;
		memory[16'h152e] <= 8'hed;
		memory[16'h152f] <= 8'hc;
		memory[16'h1530] <= 8'h5;
		memory[16'h1531] <= 8'hbc;
		memory[16'h1532] <= 8'hb3;
		memory[16'h1533] <= 8'h3e;
		memory[16'h1534] <= 8'h24;
		memory[16'h1535] <= 8'h0;
		memory[16'h1536] <= 8'ha0;
		memory[16'h1537] <= 8'h4a;
		memory[16'h1538] <= 8'h97;
		memory[16'h1539] <= 8'h39;
		memory[16'h153a] <= 8'h7b;
		memory[16'h153b] <= 8'h74;
		memory[16'h153c] <= 8'h63;
		memory[16'h153d] <= 8'hb0;
		memory[16'h153e] <= 8'hbe;
		memory[16'h153f] <= 8'h90;
		memory[16'h1540] <= 8'hc3;
		memory[16'h1541] <= 8'h1c;
		memory[16'h1542] <= 8'h62;
		memory[16'h1543] <= 8'hd7;
		memory[16'h1544] <= 8'h59;
		memory[16'h1545] <= 8'he9;
		memory[16'h1546] <= 8'hc3;
		memory[16'h1547] <= 8'h14;
		memory[16'h1548] <= 8'h66;
		memory[16'h1549] <= 8'h45;
		memory[16'h154a] <= 8'h4a;
		memory[16'h154b] <= 8'h80;
		memory[16'h154c] <= 8'h4c;
		memory[16'h154d] <= 8'h37;
		memory[16'h154e] <= 8'h8c;
		memory[16'h154f] <= 8'h51;
		memory[16'h1550] <= 8'hf4;
		memory[16'h1551] <= 8'h40;
		memory[16'h1552] <= 8'h8f;
		memory[16'h1553] <= 8'h18;
		memory[16'h1554] <= 8'h40;
		memory[16'h1555] <= 8'h2f;
		memory[16'h1556] <= 8'h62;
		memory[16'h1557] <= 8'hd8;
		memory[16'h1558] <= 8'h68;
		memory[16'h1559] <= 8'hdd;
		memory[16'h155a] <= 8'h4c;
		memory[16'h155b] <= 8'hcb;
		memory[16'h155c] <= 8'h8d;
		memory[16'h155d] <= 8'hb;
		memory[16'h155e] <= 8'h5c;
		memory[16'h155f] <= 8'h50;
		memory[16'h1560] <= 8'h27;
		memory[16'h1561] <= 8'hbe;
		memory[16'h1562] <= 8'h27;
		memory[16'h1563] <= 8'h80;
		memory[16'h1564] <= 8'ha7;
		memory[16'h1565] <= 8'heb;
		memory[16'h1566] <= 8'h94;
		memory[16'h1567] <= 8'he;
		memory[16'h1568] <= 8'h30;
		memory[16'h1569] <= 8'hde;
		memory[16'h156a] <= 8'h8e;
		memory[16'h156b] <= 8'h7c;
		memory[16'h156c] <= 8'h16;
		memory[16'h156d] <= 8'h1b;
		memory[16'h156e] <= 8'hcd;
		memory[16'h156f] <= 8'ha;
		memory[16'h1570] <= 8'h5b;
		memory[16'h1571] <= 8'h5d;
		memory[16'h1572] <= 8'h22;
		memory[16'h1573] <= 8'h9b;
		memory[16'h1574] <= 8'h8c;
		memory[16'h1575] <= 8'h84;
		memory[16'h1576] <= 8'h73;
		memory[16'h1577] <= 8'hf5;
		memory[16'h1578] <= 8'h62;
		memory[16'h1579] <= 8'hc0;
		memory[16'h157a] <= 8'hc0;
		memory[16'h157b] <= 8'hef;
		memory[16'h157c] <= 8'hcb;
		memory[16'h157d] <= 8'h1c;
		memory[16'h157e] <= 8'h40;
		memory[16'h157f] <= 8'hf2;
		memory[16'h1580] <= 8'hdb;
		memory[16'h1581] <= 8'h67;
		memory[16'h1582] <= 8'h73;
		memory[16'h1583] <= 8'h82;
		memory[16'h1584] <= 8'h52;
		memory[16'h1585] <= 8'h7;
		memory[16'h1586] <= 8'h90;
		memory[16'h1587] <= 8'h82;
		memory[16'h1588] <= 8'he6;
		memory[16'h1589] <= 8'h1f;
		memory[16'h158a] <= 8'hfe;
		memory[16'h158b] <= 8'hfc;
		memory[16'h158c] <= 8'h3a;
		memory[16'h158d] <= 8'hcc;
		memory[16'h158e] <= 8'h6;
		memory[16'h158f] <= 8'h95;
		memory[16'h1590] <= 8'h29;
		memory[16'h1591] <= 8'h28;
		memory[16'h1592] <= 8'h30;
		memory[16'h1593] <= 8'hb5;
		memory[16'h1594] <= 8'hac;
		memory[16'h1595] <= 8'ha4;
		memory[16'h1596] <= 8'haa;
		memory[16'h1597] <= 8'he;
		memory[16'h1598] <= 8'h64;
		memory[16'h1599] <= 8'h6b;
		memory[16'h159a] <= 8'hfe;
		memory[16'h159b] <= 8'h2f;
		memory[16'h159c] <= 8'h87;
		memory[16'h159d] <= 8'h3e;
		memory[16'h159e] <= 8'h21;
		memory[16'h159f] <= 8'h62;
		memory[16'h15a0] <= 8'ha5;
		memory[16'h15a1] <= 8'h94;
		memory[16'h15a2] <= 8'he5;
		memory[16'h15a3] <= 8'hf8;
		memory[16'h15a4] <= 8'h9c;
		memory[16'h15a5] <= 8'h75;
		memory[16'h15a6] <= 8'h7a;
		memory[16'h15a7] <= 8'h82;
		memory[16'h15a8] <= 8'h94;
		memory[16'h15a9] <= 8'h79;
		memory[16'h15aa] <= 8'h7e;
		memory[16'h15ab] <= 8'hce;
		memory[16'h15ac] <= 8'h45;
		memory[16'h15ad] <= 8'h84;
		memory[16'h15ae] <= 8'h63;
		memory[16'h15af] <= 8'h6e;
		memory[16'h15b0] <= 8'hac;
		memory[16'h15b1] <= 8'h94;
		memory[16'h15b2] <= 8'h23;
		memory[16'h15b3] <= 8'h58;
		memory[16'h15b4] <= 8'h38;
		memory[16'h15b5] <= 8'hce;
		memory[16'h15b6] <= 8'h67;
		memory[16'h15b7] <= 8'h9c;
		memory[16'h15b8] <= 8'h39;
		memory[16'h15b9] <= 8'h65;
		memory[16'h15ba] <= 8'hcb;
		memory[16'h15bb] <= 8'hc0;
		memory[16'h15bc] <= 8'ha3;
		memory[16'h15bd] <= 8'hec;
		memory[16'h15be] <= 8'h23;
		memory[16'h15bf] <= 8'h48;
		memory[16'h15c0] <= 8'h81;
		memory[16'h15c1] <= 8'h8;
		memory[16'h15c2] <= 8'h40;
		memory[16'h15c3] <= 8'h1d;
		memory[16'h15c4] <= 8'h7d;
		memory[16'h15c5] <= 8'hbb;
		memory[16'h15c6] <= 8'h9f;
		memory[16'h15c7] <= 8'h12;
		memory[16'h15c8] <= 8'h34;
		memory[16'h15c9] <= 8'h1d;
		memory[16'h15ca] <= 8'he0;
		memory[16'h15cb] <= 8'h79;
		memory[16'h15cc] <= 8'ha1;
		memory[16'h15cd] <= 8'h44;
		memory[16'h15ce] <= 8'he7;
		memory[16'h15cf] <= 8'h4d;
		memory[16'h15d0] <= 8'hd8;
		memory[16'h15d1] <= 8'ha;
		memory[16'h15d2] <= 8'ha5;
		memory[16'h15d3] <= 8'h10;
		memory[16'h15d4] <= 8'hd8;
		memory[16'h15d5] <= 8'hc;
		memory[16'h15d6] <= 8'hac;
		memory[16'h15d7] <= 8'h11;
		memory[16'h15d8] <= 8'h71;
		memory[16'h15d9] <= 8'h77;
		memory[16'h15da] <= 8'hd2;
		memory[16'h15db] <= 8'h14;
		memory[16'h15dc] <= 8'h63;
		memory[16'h15dd] <= 8'hf5;
		memory[16'h15de] <= 8'h5d;
		memory[16'h15df] <= 8'he4;
		memory[16'h15e0] <= 8'hfd;
		memory[16'h15e1] <= 8'h9d;
		memory[16'h15e2] <= 8'h1;
		memory[16'h15e3] <= 8'h7a;
		memory[16'h15e4] <= 8'h58;
		memory[16'h15e5] <= 8'ha0;
		memory[16'h15e6] <= 8'h8c;
		memory[16'h15e7] <= 8'h8c;
		memory[16'h15e8] <= 8'hbd;
		memory[16'h15e9] <= 8'h6d;
		memory[16'h15ea] <= 8'h5;
		memory[16'h15eb] <= 8'h5e;
		memory[16'h15ec] <= 8'hb1;
		memory[16'h15ed] <= 8'hec;
		memory[16'h15ee] <= 8'hab;
		memory[16'h15ef] <= 8'h89;
		memory[16'h15f0] <= 8'hf7;
		memory[16'h15f1] <= 8'h51;
		memory[16'h15f2] <= 8'h99;
		memory[16'h15f3] <= 8'hcf;
		memory[16'h15f4] <= 8'h5d;
		memory[16'h15f5] <= 8'h45;
		memory[16'h15f6] <= 8'he1;
		memory[16'h15f7] <= 8'hcf;
		memory[16'h15f8] <= 8'hbc;
		memory[16'h15f9] <= 8'hb3;
		memory[16'h15fa] <= 8'he3;
		memory[16'h15fb] <= 8'h1f;
		memory[16'h15fc] <= 8'ha8;
		memory[16'h15fd] <= 8'h40;
		memory[16'h15fe] <= 8'h4;
		memory[16'h15ff] <= 8'ha5;
		memory[16'h1600] <= 8'hde;
		memory[16'h1601] <= 8'h5;
		memory[16'h1602] <= 8'h1f;
		memory[16'h1603] <= 8'h36;
		memory[16'h1604] <= 8'ha6;
		memory[16'h1605] <= 8'hac;
		memory[16'h1606] <= 8'hc3;
		memory[16'h1607] <= 8'h63;
		memory[16'h1608] <= 8'h19;
		memory[16'h1609] <= 8'hc8;
		memory[16'h160a] <= 8'hc2;
		memory[16'h160b] <= 8'hca;
		memory[16'h160c] <= 8'hb5;
		memory[16'h160d] <= 8'h6d;
		memory[16'h160e] <= 8'h53;
		memory[16'h160f] <= 8'hac;
		memory[16'h1610] <= 8'hbe;
		memory[16'h1611] <= 8'hec;
		memory[16'h1612] <= 8'h7b;
		memory[16'h1613] <= 8'h1c;
		memory[16'h1614] <= 8'h31;
		memory[16'h1615] <= 8'h5c;
		memory[16'h1616] <= 8'heb;
		memory[16'h1617] <= 8'hed;
		memory[16'h1618] <= 8'hf;
		memory[16'h1619] <= 8'hce;
		memory[16'h161a] <= 8'hc;
		memory[16'h161b] <= 8'hb7;
		memory[16'h161c] <= 8'hf;
		memory[16'h161d] <= 8'h10;
		memory[16'h161e] <= 8'h5c;
		memory[16'h161f] <= 8'hed;
		memory[16'h1620] <= 8'h16;
		memory[16'h1621] <= 8'h7c;
		memory[16'h1622] <= 8'h23;
		memory[16'h1623] <= 8'hbc;
		memory[16'h1624] <= 8'h28;
		memory[16'h1625] <= 8'he6;
		memory[16'h1626] <= 8'h1f;
		memory[16'h1627] <= 8'h41;
		memory[16'h1628] <= 8'haf;
		memory[16'h1629] <= 8'he1;
		memory[16'h162a] <= 8'hb;
		memory[16'h162b] <= 8'h64;
		memory[16'h162c] <= 8'h4f;
		memory[16'h162d] <= 8'h5e;
		memory[16'h162e] <= 8'h10;
		memory[16'h162f] <= 8'hd;
		memory[16'h1630] <= 8'h4a;
		memory[16'h1631] <= 8'h8b;
		memory[16'h1632] <= 8'h29;
		memory[16'h1633] <= 8'h7b;
		memory[16'h1634] <= 8'he8;
		memory[16'h1635] <= 8'h14;
		memory[16'h1636] <= 8'h68;
		memory[16'h1637] <= 8'hf7;
		memory[16'h1638] <= 8'he3;
		memory[16'h1639] <= 8'h74;
		memory[16'h163a] <= 8'haf;
		memory[16'h163b] <= 8'hf2;
		memory[16'h163c] <= 8'h85;
		memory[16'h163d] <= 8'hb;
		memory[16'h163e] <= 8'hdf;
		memory[16'h163f] <= 8'h9b;
		memory[16'h1640] <= 8'h87;
		memory[16'h1641] <= 8'h2;
		memory[16'h1642] <= 8'h57;
		memory[16'h1643] <= 8'haf;
		memory[16'h1644] <= 8'he9;
		memory[16'h1645] <= 8'h76;
		memory[16'h1646] <= 8'hf0;
		memory[16'h1647] <= 8'h98;
		memory[16'h1648] <= 8'h58;
		memory[16'h1649] <= 8'hfb;
		memory[16'h164a] <= 8'hfc;
		memory[16'h164b] <= 8'ha7;
		memory[16'h164c] <= 8'h59;
		memory[16'h164d] <= 8'hc;
		memory[16'h164e] <= 8'hb4;
		memory[16'h164f] <= 8'ha3;
		memory[16'h1650] <= 8'h97;
		memory[16'h1651] <= 8'hde;
		memory[16'h1652] <= 8'h1e;
		memory[16'h1653] <= 8'h7f;
		memory[16'h1654] <= 8'hf2;
		memory[16'h1655] <= 8'h86;
		memory[16'h1656] <= 8'h77;
		memory[16'h1657] <= 8'hd5;
		memory[16'h1658] <= 8'hfb;
		memory[16'h1659] <= 8'h26;
		memory[16'h165a] <= 8'hc7;
		memory[16'h165b] <= 8'h80;
		memory[16'h165c] <= 8'h31;
		memory[16'h165d] <= 8'ha6;
		memory[16'h165e] <= 8'h1b;
		memory[16'h165f] <= 8'hb9;
		memory[16'h1660] <= 8'ha9;
		memory[16'h1661] <= 8'h72;
		memory[16'h1662] <= 8'h68;
		memory[16'h1663] <= 8'h92;
		memory[16'h1664] <= 8'he8;
		memory[16'h1665] <= 8'h59;
		memory[16'h1666] <= 8'h2a;
		memory[16'h1667] <= 8'h40;
		memory[16'h1668] <= 8'h54;
		memory[16'h1669] <= 8'h26;
		memory[16'h166a] <= 8'he7;
		memory[16'h166b] <= 8'hae;
		memory[16'h166c] <= 8'h32;
		memory[16'h166d] <= 8'h9c;
		memory[16'h166e] <= 8'h51;
		memory[16'h166f] <= 8'hc9;
		memory[16'h1670] <= 8'h7a;
		memory[16'h1671] <= 8'h70;
		memory[16'h1672] <= 8'h49;
		memory[16'h1673] <= 8'h6c;
		memory[16'h1674] <= 8'hf6;
		memory[16'h1675] <= 8'hc0;
		memory[16'h1676] <= 8'h42;
		memory[16'h1677] <= 8'hf1;
		memory[16'h1678] <= 8'he6;
		memory[16'h1679] <= 8'h9;
		memory[16'h167a] <= 8'h71;
		memory[16'h167b] <= 8'h17;
		memory[16'h167c] <= 8'hb0;
		memory[16'h167d] <= 8'h8c;
		memory[16'h167e] <= 8'hd0;
		memory[16'h167f] <= 8'h59;
		memory[16'h1680] <= 8'hfe;
		memory[16'h1681] <= 8'h39;
		memory[16'h1682] <= 8'heb;
		memory[16'h1683] <= 8'he7;
		memory[16'h1684] <= 8'h92;
		memory[16'h1685] <= 8'h15;
		memory[16'h1686] <= 8'h27;
		memory[16'h1687] <= 8'he6;
		memory[16'h1688] <= 8'h3b;
		memory[16'h1689] <= 8'hf;
		memory[16'h168a] <= 8'h94;
		memory[16'h168b] <= 8'h6d;
		memory[16'h168c] <= 8'hab;
		memory[16'h168d] <= 8'he6;
		memory[16'h168e] <= 8'h36;
		memory[16'h168f] <= 8'h25;
		memory[16'h1690] <= 8'h56;
		memory[16'h1691] <= 8'h7f;
		memory[16'h1692] <= 8'h91;
		memory[16'h1693] <= 8'h4c;
		memory[16'h1694] <= 8'h3f;
		memory[16'h1695] <= 8'hd3;
		memory[16'h1696] <= 8'h3e;
		memory[16'h1697] <= 8'h25;
		memory[16'h1698] <= 8'hdd;
		memory[16'h1699] <= 8'haf;
		memory[16'h169a] <= 8'h3d;
		memory[16'h169b] <= 8'h8d;
		memory[16'h169c] <= 8'h3c;
		memory[16'h169d] <= 8'hd;
		memory[16'h169e] <= 8'he6;
		memory[16'h169f] <= 8'h3a;
		memory[16'h16a0] <= 8'h46;
		memory[16'h16a1] <= 8'hd1;
		memory[16'h16a2] <= 8'h21;
		memory[16'h16a3] <= 8'hd8;
		memory[16'h16a4] <= 8'he6;
		memory[16'h16a5] <= 8'h49;
		memory[16'h16a6] <= 8'hbf;
		memory[16'h16a7] <= 8'h21;
		memory[16'h16a8] <= 8'h58;
		memory[16'h16a9] <= 8'h53;
		memory[16'h16aa] <= 8'h8e;
		memory[16'h16ab] <= 8'h3;
		memory[16'h16ac] <= 8'h39;
		memory[16'h16ad] <= 8'hc4;
		memory[16'h16ae] <= 8'h28;
		memory[16'h16af] <= 8'h8f;
		memory[16'h16b0] <= 8'h44;
		memory[16'h16b1] <= 8'hb9;
		memory[16'h16b2] <= 8'hdc;
		memory[16'h16b3] <= 8'h83;
		memory[16'h16b4] <= 8'h8d;
		memory[16'h16b5] <= 8'h1a;
		memory[16'h16b6] <= 8'ha9;
		memory[16'h16b7] <= 8'h6a;
		memory[16'h16b8] <= 8'hc9;
		memory[16'h16b9] <= 8'he6;
		memory[16'h16ba] <= 8'hf7;
		memory[16'h16bb] <= 8'h5;
		memory[16'h16bc] <= 8'hf3;
		memory[16'h16bd] <= 8'hdd;
		memory[16'h16be] <= 8'h40;
		memory[16'h16bf] <= 8'h3a;
		memory[16'h16c0] <= 8'hae;
		memory[16'h16c1] <= 8'h61;
		memory[16'h16c2] <= 8'h12;
		memory[16'h16c3] <= 8'h94;
		memory[16'h16c4] <= 8'haa;
		memory[16'h16c5] <= 8'hd1;
		memory[16'h16c6] <= 8'hb5;
		memory[16'h16c7] <= 8'h2;
		memory[16'h16c8] <= 8'h25;
		memory[16'h16c9] <= 8'h43;
		memory[16'h16ca] <= 8'h5;
		memory[16'h16cb] <= 8'h5e;
		memory[16'h16cc] <= 8'h7;
		memory[16'h16cd] <= 8'h2d;
		memory[16'h16ce] <= 8'hee;
		memory[16'h16cf] <= 8'h4b;
		memory[16'h16d0] <= 8'he7;
		memory[16'h16d1] <= 8'hca;
		memory[16'h16d2] <= 8'hcf;
		memory[16'h16d3] <= 8'h74;
		memory[16'h16d4] <= 8'he4;
		memory[16'h16d5] <= 8'h78;
		memory[16'h16d6] <= 8'hde;
		memory[16'h16d7] <= 8'had;
		memory[16'h16d8] <= 8'h5e;
		memory[16'h16d9] <= 8'hd5;
		memory[16'h16da] <= 8'hb3;
		memory[16'h16db] <= 8'h51;
		memory[16'h16dc] <= 8'hb2;
		memory[16'h16dd] <= 8'hf3;
		memory[16'h16de] <= 8'h8b;
		memory[16'h16df] <= 8'h60;
		memory[16'h16e0] <= 8'h54;
		memory[16'h16e1] <= 8'h9e;
		memory[16'h16e2] <= 8'hf4;
		memory[16'h16e3] <= 8'hff;
		memory[16'h16e4] <= 8'h6f;
		memory[16'h16e5] <= 8'ha9;
		memory[16'h16e6] <= 8'h1;
		memory[16'h16e7] <= 8'h94;
		memory[16'h16e8] <= 8'hec;
		memory[16'h16e9] <= 8'h7;
		memory[16'h16ea] <= 8'hf3;
		memory[16'h16eb] <= 8'hf3;
		memory[16'h16ec] <= 8'h34;
		memory[16'h16ed] <= 8'he1;
		memory[16'h16ee] <= 8'h3f;
		memory[16'h16ef] <= 8'h1b;
		memory[16'h16f0] <= 8'hab;
		memory[16'h16f1] <= 8'he;
		memory[16'h16f2] <= 8'h8f;
		memory[16'h16f3] <= 8'h8f;
		memory[16'h16f4] <= 8'h86;
		memory[16'h16f5] <= 8'h6d;
		memory[16'h16f6] <= 8'h3c;
		memory[16'h16f7] <= 8'he4;
		memory[16'h16f8] <= 8'h42;
		memory[16'h16f9] <= 8'hef;
		memory[16'h16fa] <= 8'h35;
		memory[16'h16fb] <= 8'hf4;
		memory[16'h16fc] <= 8'he2;
		memory[16'h16fd] <= 8'hc1;
		memory[16'h16fe] <= 8'h54;
		memory[16'h16ff] <= 8'h37;
		memory[16'h1700] <= 8'h5f;
		memory[16'h1701] <= 8'h48;
		memory[16'h1702] <= 8'h36;
		memory[16'h1703] <= 8'hce;
		memory[16'h1704] <= 8'hf1;
		memory[16'h1705] <= 8'h37;
		memory[16'h1706] <= 8'h63;
		memory[16'h1707] <= 8'hdd;
		memory[16'h1708] <= 8'h3e;
		memory[16'h1709] <= 8'h56;
		memory[16'h170a] <= 8'hd1;
		memory[16'h170b] <= 8'h73;
		memory[16'h170c] <= 8'h37;
		memory[16'h170d] <= 8'h10;
		memory[16'h170e] <= 8'h8e;
		memory[16'h170f] <= 8'he2;
		memory[16'h1710] <= 8'h1e;
		memory[16'h1711] <= 8'h1e;
		memory[16'h1712] <= 8'h71;
		memory[16'h1713] <= 8'ha4;
		memory[16'h1714] <= 8'h8b;
		memory[16'h1715] <= 8'had;
		memory[16'h1716] <= 8'h88;
		memory[16'h1717] <= 8'hce;
		memory[16'h1718] <= 8'h9d;
		memory[16'h1719] <= 8'hbd;
		memory[16'h171a] <= 8'hc2;
		memory[16'h171b] <= 8'h7f;
		memory[16'h171c] <= 8'h7e;
		memory[16'h171d] <= 8'h17;
		memory[16'h171e] <= 8'hb6;
		memory[16'h171f] <= 8'hdd;
		memory[16'h1720] <= 8'h5f;
		memory[16'h1721] <= 8'hec;
		memory[16'h1722] <= 8'hac;
		memory[16'h1723] <= 8'h51;
		memory[16'h1724] <= 8'h24;
		memory[16'h1725] <= 8'hf;
		memory[16'h1726] <= 8'h2e;
		memory[16'h1727] <= 8'h62;
		memory[16'h1728] <= 8'h65;
		memory[16'h1729] <= 8'hff;
		memory[16'h172a] <= 8'hd5;
		memory[16'h172b] <= 8'h9c;
		memory[16'h172c] <= 8'hf;
		memory[16'h172d] <= 8'h64;
		memory[16'h172e] <= 8'h7e;
		memory[16'h172f] <= 8'h2d;
		memory[16'h1730] <= 8'h82;
		memory[16'h1731] <= 8'hef;
		memory[16'h1732] <= 8'hd1;
		memory[16'h1733] <= 8'hd;
		memory[16'h1734] <= 8'h9c;
		memory[16'h1735] <= 8'h59;
		memory[16'h1736] <= 8'hdb;
		memory[16'h1737] <= 8'h39;
		memory[16'h1738] <= 8'h17;
		memory[16'h1739] <= 8'h9e;
		memory[16'h173a] <= 8'hb9;
		memory[16'h173b] <= 8'h95;
		memory[16'h173c] <= 8'hb5;
		memory[16'h173d] <= 8'h6f;
		memory[16'h173e] <= 8'h73;
		memory[16'h173f] <= 8'h14;
		memory[16'h1740] <= 8'h5c;
		memory[16'h1741] <= 8'h1f;
		memory[16'h1742] <= 8'h65;
		memory[16'h1743] <= 8'h80;
		memory[16'h1744] <= 8'h2e;
		memory[16'h1745] <= 8'h94;
		memory[16'h1746] <= 8'he2;
		memory[16'h1747] <= 8'h93;
		memory[16'h1748] <= 8'h93;
		memory[16'h1749] <= 8'hb8;
		memory[16'h174a] <= 8'h2f;
		memory[16'h174b] <= 8'ha3;
		memory[16'h174c] <= 8'h1c;
		memory[16'h174d] <= 8'had;
		memory[16'h174e] <= 8'hd0;
		memory[16'h174f] <= 8'h9e;
		memory[16'h1750] <= 8'h9c;
		memory[16'h1751] <= 8'ha2;
		memory[16'h1752] <= 8'hab;
		memory[16'h1753] <= 8'h38;
		memory[16'h1754] <= 8'hfb;
		memory[16'h1755] <= 8'h87;
		memory[16'h1756] <= 8'h72;
		memory[16'h1757] <= 8'h12;
		memory[16'h1758] <= 8'h25;
		memory[16'h1759] <= 8'h2b;
		memory[16'h175a] <= 8'ha8;
		memory[16'h175b] <= 8'hda;
		memory[16'h175c] <= 8'h9a;
		memory[16'h175d] <= 8'h1b;
		memory[16'h175e] <= 8'hee;
		memory[16'h175f] <= 8'hf6;
		memory[16'h1760] <= 8'h3a;
		memory[16'h1761] <= 8'h54;
		memory[16'h1762] <= 8'h76;
		memory[16'h1763] <= 8'h68;
		memory[16'h1764] <= 8'he8;
		memory[16'h1765] <= 8'h59;
		memory[16'h1766] <= 8'hfb;
		memory[16'h1767] <= 8'h7b;
		memory[16'h1768] <= 8'h11;
		memory[16'h1769] <= 8'h2a;
		memory[16'h176a] <= 8'h1e;
		memory[16'h176b] <= 8'h2d;
		memory[16'h176c] <= 8'hd7;
		memory[16'h176d] <= 8'hef;
		memory[16'h176e] <= 8'hcb;
		memory[16'h176f] <= 8'h73;
		memory[16'h1770] <= 8'h91;
		memory[16'h1771] <= 8'h76;
		memory[16'h1772] <= 8'hab;
		memory[16'h1773] <= 8'h8c;
		memory[16'h1774] <= 8'hfd;
		memory[16'h1775] <= 8'h1d;
		memory[16'h1776] <= 8'h9f;
		memory[16'h1777] <= 8'h22;
		memory[16'h1778] <= 8'h48;
		memory[16'h1779] <= 8'h47;
		memory[16'h177a] <= 8'hfc;
		memory[16'h177b] <= 8'he3;
		memory[16'h177c] <= 8'h62;
		memory[16'h177d] <= 8'heb;
		memory[16'h177e] <= 8'hd9;
		memory[16'h177f] <= 8'h9c;
		memory[16'h1780] <= 8'h3f;
		memory[16'h1781] <= 8'h50;
		memory[16'h1782] <= 8'h4;
		memory[16'h1783] <= 8'h27;
		memory[16'h1784] <= 8'ha9;
		memory[16'h1785] <= 8'hff;
		memory[16'h1786] <= 8'ha2;
		memory[16'h1787] <= 8'hba;
		memory[16'h1788] <= 8'h29;
		memory[16'h1789] <= 8'hc1;
		memory[16'h178a] <= 8'he7;
		memory[16'h178b] <= 8'h0;
		memory[16'h178c] <= 8'hb0;
		memory[16'h178d] <= 8'hb2;
		memory[16'h178e] <= 8'h73;
		memory[16'h178f] <= 8'h41;
		memory[16'h1790] <= 8'h28;
		memory[16'h1791] <= 8'h1e;
		memory[16'h1792] <= 8'hcd;
		memory[16'h1793] <= 8'h26;
		memory[16'h1794] <= 8'h3c;
		memory[16'h1795] <= 8'h6c;
		memory[16'h1796] <= 8'h48;
		memory[16'h1797] <= 8'h84;
		memory[16'h1798] <= 8'hb3;
		memory[16'h1799] <= 8'h45;
		memory[16'h179a] <= 8'h67;
		memory[16'h179b] <= 8'h15;
		memory[16'h179c] <= 8'h30;
		memory[16'h179d] <= 8'h41;
		memory[16'h179e] <= 8'hb1;
		memory[16'h179f] <= 8'h6f;
		memory[16'h17a0] <= 8'h91;
		memory[16'h17a1] <= 8'hb5;
		memory[16'h17a2] <= 8'h96;
		memory[16'h17a3] <= 8'h3a;
		memory[16'h17a4] <= 8'hb4;
		memory[16'h17a5] <= 8'h38;
		memory[16'h17a6] <= 8'hf4;
		memory[16'h17a7] <= 8'hdd;
		memory[16'h17a8] <= 8'hf9;
		memory[16'h17a9] <= 8'hdb;
		memory[16'h17aa] <= 8'hdd;
		memory[16'h17ab] <= 8'ha9;
		memory[16'h17ac] <= 8'h8d;
		memory[16'h17ad] <= 8'h50;
		memory[16'h17ae] <= 8'hea;
		memory[16'h17af] <= 8'hb5;
		memory[16'h17b0] <= 8'h6f;
		memory[16'h17b1] <= 8'hb8;
		memory[16'h17b2] <= 8'hdb;
		memory[16'h17b3] <= 8'hab;
		memory[16'h17b4] <= 8'h24;
		memory[16'h17b5] <= 8'h24;
		memory[16'h17b6] <= 8'h2f;
		memory[16'h17b7] <= 8'hd8;
		memory[16'h17b8] <= 8'h69;
		memory[16'h17b9] <= 8'h97;
		memory[16'h17ba] <= 8'hed;
		memory[16'h17bb] <= 8'h99;
		memory[16'h17bc] <= 8'hd8;
		memory[16'h17bd] <= 8'h9f;
		memory[16'h17be] <= 8'h8;
		memory[16'h17bf] <= 8'h69;
		memory[16'h17c0] <= 8'h54;
		memory[16'h17c1] <= 8'h9e;
		memory[16'h17c2] <= 8'ha3;
		memory[16'h17c3] <= 8'h9;
		memory[16'h17c4] <= 8'hd6;
		memory[16'h17c5] <= 8'h97;
		memory[16'h17c6] <= 8'he6;
		memory[16'h17c7] <= 8'hd0;
		memory[16'h17c8] <= 8'h72;
		memory[16'h17c9] <= 8'hc4;
		memory[16'h17ca] <= 8'h79;
		memory[16'h17cb] <= 8'hff;
		memory[16'h17cc] <= 8'h14;
		memory[16'h17cd] <= 8'h64;
		memory[16'h17ce] <= 8'hb4;
		memory[16'h17cf] <= 8'h83;
		memory[16'h17d0] <= 8'h1c;
		memory[16'h17d1] <= 8'h90;
		memory[16'h17d2] <= 8'h2e;
		memory[16'h17d3] <= 8'h40;
		memory[16'h17d4] <= 8'hb4;
		memory[16'h17d5] <= 8'h5e;
		memory[16'h17d6] <= 8'h18;
		memory[16'h17d7] <= 8'h1d;
		memory[16'h17d8] <= 8'hf5;
		memory[16'h17d9] <= 8'h6;
		memory[16'h17da] <= 8'hb6;
		memory[16'h17db] <= 8'hcd;
		memory[16'h17dc] <= 8'ha5;
		memory[16'h17dd] <= 8'hbe;
		memory[16'h17de] <= 8'h36;
		memory[16'h17df] <= 8'hf9;
		memory[16'h17e0] <= 8'h5c;
		memory[16'h17e1] <= 8'hd9;
		memory[16'h17e2] <= 8'h2;
		memory[16'h17e3] <= 8'h32;
		memory[16'h17e4] <= 8'h70;
		memory[16'h17e5] <= 8'he9;
		memory[16'h17e6] <= 8'h2;
		memory[16'h17e7] <= 8'he2;
		memory[16'h17e8] <= 8'had;
		memory[16'h17e9] <= 8'h7c;
		memory[16'h17ea] <= 8'he1;
		memory[16'h17eb] <= 8'hc1;
		memory[16'h17ec] <= 8'he0;
		memory[16'h17ed] <= 8'h95;
		memory[16'h17ee] <= 8'h45;
		memory[16'h17ef] <= 8'hfc;
		memory[16'h17f0] <= 8'h25;
		memory[16'h17f1] <= 8'h73;
		memory[16'h17f2] <= 8'h3c;
		memory[16'h17f3] <= 8'hd9;
		memory[16'h17f4] <= 8'hd1;
		memory[16'h17f5] <= 8'h55;
		memory[16'h17f6] <= 8'hf6;
		memory[16'h17f7] <= 8'hc6;
		memory[16'h17f8] <= 8'h5b;
		memory[16'h17f9] <= 8'hac;
		memory[16'h17fa] <= 8'h93;
		memory[16'h17fb] <= 8'h0;
		memory[16'h17fc] <= 8'h6a;
		memory[16'h17fd] <= 8'hc9;
		memory[16'h17fe] <= 8'hf9;
		memory[16'h17ff] <= 8'hc6;
		memory[16'h1800] <= 8'ha2;
		memory[16'h1801] <= 8'hfc;
		memory[16'h1802] <= 8'hf9;
		memory[16'h1803] <= 8'h12;
		memory[16'h1804] <= 8'he5;
		memory[16'h1805] <= 8'hfb;
		memory[16'h1806] <= 8'hf4;
		memory[16'h1807] <= 8'h92;
		memory[16'h1808] <= 8'h77;
		memory[16'h1809] <= 8'hd5;
		memory[16'h180a] <= 8'h53;
		memory[16'h180b] <= 8'h57;
		memory[16'h180c] <= 8'h6b;
		memory[16'h180d] <= 8'h98;
		memory[16'h180e] <= 8'h53;
		memory[16'h180f] <= 8'h90;
		memory[16'h1810] <= 8'hc;
		memory[16'h1811] <= 8'h90;
		memory[16'h1812] <= 8'h6a;
		memory[16'h1813] <= 8'hdd;
		memory[16'h1814] <= 8'he5;
		memory[16'h1815] <= 8'h60;
		memory[16'h1816] <= 8'ha4;
		memory[16'h1817] <= 8'h40;
		memory[16'h1818] <= 8'hd;
		memory[16'h1819] <= 8'h37;
		memory[16'h181a] <= 8'h40;
		memory[16'h181b] <= 8'h77;
		memory[16'h181c] <= 8'h1;
		memory[16'h181d] <= 8'h39;
		memory[16'h181e] <= 8'h3e;
		memory[16'h181f] <= 8'ha3;
		memory[16'h1820] <= 8'h35;
		memory[16'h1821] <= 8'h37;
		memory[16'h1822] <= 8'hb6;
		memory[16'h1823] <= 8'h1a;
		memory[16'h1824] <= 8'h32;
		memory[16'h1825] <= 8'haa;
		memory[16'h1826] <= 8'hac;
		memory[16'h1827] <= 8'haa;
		memory[16'h1828] <= 8'h80;
		memory[16'h1829] <= 8'h0;
		memory[16'h182a] <= 8'h1;
		memory[16'h182b] <= 8'heb;
		memory[16'h182c] <= 8'h98;
		memory[16'h182d] <= 8'h55;
		memory[16'h182e] <= 8'h7b;
		memory[16'h182f] <= 8'ha4;
		memory[16'h1830] <= 8'he5;
		memory[16'h1831] <= 8'he5;
		memory[16'h1832] <= 8'h82;
		memory[16'h1833] <= 8'hca;
		memory[16'h1834] <= 8'h46;
		memory[16'h1835] <= 8'h26;
		memory[16'h1836] <= 8'ha;
		memory[16'h1837] <= 8'h53;
		memory[16'h1838] <= 8'h5d;
		memory[16'h1839] <= 8'h4a;
		memory[16'h183a] <= 8'hca;
		memory[16'h183b] <= 8'h5e;
		memory[16'h183c] <= 8'h83;
		memory[16'h183d] <= 8'h8;
		memory[16'h183e] <= 8'h2;
		memory[16'h183f] <= 8'hb9;
		memory[16'h1840] <= 8'h3f;
		memory[16'h1841] <= 8'hb8;
		memory[16'h1842] <= 8'hd3;
		memory[16'h1843] <= 8'h72;
		memory[16'h1844] <= 8'h62;
		memory[16'h1845] <= 8'h80;
		memory[16'h1846] <= 8'h1c;
		memory[16'h1847] <= 8'he2;
		memory[16'h1848] <= 8'h80;
		memory[16'h1849] <= 8'h1d;
		memory[16'h184a] <= 8'hcd;
		memory[16'h184b] <= 8'h18;
		memory[16'h184c] <= 8'h72;
		memory[16'h184d] <= 8'h49;
		memory[16'h184e] <= 8'hbd;
		memory[16'h184f] <= 8'h57;
		memory[16'h1850] <= 8'h2e;
		memory[16'h1851] <= 8'h3f;
		memory[16'h1852] <= 8'h21;
		memory[16'h1853] <= 8'h74;
		memory[16'h1854] <= 8'h65;
		memory[16'h1855] <= 8'h2b;
		memory[16'h1856] <= 8'hc7;
		memory[16'h1857] <= 8'hc2;
		memory[16'h1858] <= 8'h75;
		memory[16'h1859] <= 8'h92;
		memory[16'h185a] <= 8'h21;
		memory[16'h185b] <= 8'hf9;
		memory[16'h185c] <= 8'h9a;
		memory[16'h185d] <= 8'h23;
		memory[16'h185e] <= 8'hb2;
		memory[16'h185f] <= 8'hda;
		memory[16'h1860] <= 8'hdb;
		memory[16'h1861] <= 8'h85;
		memory[16'h1862] <= 8'h4c;
		memory[16'h1863] <= 8'h3d;
		memory[16'h1864] <= 8'h5;
		memory[16'h1865] <= 8'h68;
		memory[16'h1866] <= 8'h20;
		memory[16'h1867] <= 8'h85;
		memory[16'h1868] <= 8'h85;
		memory[16'h1869] <= 8'hed;
		memory[16'h186a] <= 8'h9e;
		memory[16'h186b] <= 8'hf8;
		memory[16'h186c] <= 8'h36;
		memory[16'h186d] <= 8'h5b;
		memory[16'h186e] <= 8'h4f;
		memory[16'h186f] <= 8'h65;
		memory[16'h1870] <= 8'h9a;
		memory[16'h1871] <= 8'h71;
		memory[16'h1872] <= 8'hd9;
		memory[16'h1873] <= 8'hff;
		memory[16'h1874] <= 8'h9c;
		memory[16'h1875] <= 8'ha1;
		memory[16'h1876] <= 8'hc1;
		memory[16'h1877] <= 8'h12;
		memory[16'h1878] <= 8'h33;
		memory[16'h1879] <= 8'he2;
		memory[16'h187a] <= 8'hb;
		memory[16'h187b] <= 8'hcd;
		memory[16'h187c] <= 8'h5;
		memory[16'h187d] <= 8'hbd;
		memory[16'h187e] <= 8'ha7;
		memory[16'h187f] <= 8'he0;
		memory[16'h1880] <= 8'h42;
		memory[16'h1881] <= 8'hf3;
		memory[16'h1882] <= 8'h1e;
		memory[16'h1883] <= 8'h48;
		memory[16'h1884] <= 8'h5b;
		memory[16'h1885] <= 8'h3e;
		memory[16'h1886] <= 8'hcd;
		memory[16'h1887] <= 8'he1;
		memory[16'h1888] <= 8'h2b;
		memory[16'h1889] <= 8'h6b;
		memory[16'h188a] <= 8'hd9;
		memory[16'h188b] <= 8'h62;
		memory[16'h188c] <= 8'hc6;
		memory[16'h188d] <= 8'h28;
		memory[16'h188e] <= 8'hc7;
		memory[16'h188f] <= 8'h60;
		memory[16'h1890] <= 8'h99;
		memory[16'h1891] <= 8'ha0;
		memory[16'h1892] <= 8'h5f;
		memory[16'h1893] <= 8'h36;
		memory[16'h1894] <= 8'h41;
		memory[16'h1895] <= 8'h21;
		memory[16'h1896] <= 8'h48;
		memory[16'h1897] <= 8'h74;
		memory[16'h1898] <= 8'h3;
		memory[16'h1899] <= 8'h53;
		memory[16'h189a] <= 8'h42;
		memory[16'h189b] <= 8'h9;
		memory[16'h189c] <= 8'h10;
		memory[16'h189d] <= 8'he9;
		memory[16'h189e] <= 8'he9;
		memory[16'h189f] <= 8'h52;
		memory[16'h18a0] <= 8'hdd;
		memory[16'h18a1] <= 8'h7;
		memory[16'h18a2] <= 8'h9a;
		memory[16'h18a3] <= 8'h38;
		memory[16'h18a4] <= 8'h45;
		memory[16'h18a5] <= 8'h68;
		memory[16'h18a6] <= 8'h19;
		memory[16'h18a7] <= 8'h71;
		memory[16'h18a8] <= 8'hd3;
		memory[16'h18a9] <= 8'hf2;
		memory[16'h18aa] <= 8'hd3;
		memory[16'h18ab] <= 8'h9a;
		memory[16'h18ac] <= 8'h1b;
		memory[16'h18ad] <= 8'h9a;
		memory[16'h18ae] <= 8'hfa;
		memory[16'h18af] <= 8'hb4;
		memory[16'h18b0] <= 8'h3a;
		memory[16'h18b1] <= 8'h5a;
		memory[16'h18b2] <= 8'hea;
		memory[16'h18b3] <= 8'h7c;
		memory[16'h18b4] <= 8'h7b;
		memory[16'h18b5] <= 8'h32;
		memory[16'h18b6] <= 8'hf0;
		memory[16'h18b7] <= 8'h7e;
		memory[16'h18b8] <= 8'h85;
		memory[16'h18b9] <= 8'h32;
		memory[16'h18ba] <= 8'h87;
		memory[16'h18bb] <= 8'h95;
		memory[16'h18bc] <= 8'h1c;
		memory[16'h18bd] <= 8'h71;
		memory[16'h18be] <= 8'he8;
		memory[16'h18bf] <= 8'hf9;
		memory[16'h18c0] <= 8'h78;
		memory[16'h18c1] <= 8'h82;
		memory[16'h18c2] <= 8'h31;
		memory[16'h18c3] <= 8'hbe;
		memory[16'h18c4] <= 8'hea;
		memory[16'h18c5] <= 8'h4b;
		memory[16'h18c6] <= 8'h2f;
		memory[16'h18c7] <= 8'hbe;
		memory[16'h18c8] <= 8'h3d;
		memory[16'h18c9] <= 8'h2;
		memory[16'h18ca] <= 8'h58;
		memory[16'h18cb] <= 8'h58;
		memory[16'h18cc] <= 8'h9c;
		memory[16'h18cd] <= 8'h52;
		memory[16'h18ce] <= 8'hd;
		memory[16'h18cf] <= 8'hd6;
		memory[16'h18d0] <= 8'hac;
		memory[16'h18d1] <= 8'hf7;
		memory[16'h18d2] <= 8'h52;
		memory[16'h18d3] <= 8'h27;
		memory[16'h18d4] <= 8'h2a;
		memory[16'h18d5] <= 8'h43;
		memory[16'h18d6] <= 8'ha6;
		memory[16'h18d7] <= 8'haf;
		memory[16'h18d8] <= 8'h75;
		memory[16'h18d9] <= 8'h2d;
		memory[16'h18da] <= 8'h45;
		memory[16'h18db] <= 8'h91;
		memory[16'h18dc] <= 8'h9e;
		memory[16'h18dd] <= 8'h2d;
		memory[16'h18de] <= 8'h8a;
		memory[16'h18df] <= 8'h17;
		memory[16'h18e0] <= 8'haf;
		memory[16'h18e1] <= 8'hbc;
		memory[16'h18e2] <= 8'hd5;
		memory[16'h18e3] <= 8'h9a;
		memory[16'h18e4] <= 8'h7;
		memory[16'h18e5] <= 8'h4;
		memory[16'h18e6] <= 8'h58;
		memory[16'h18e7] <= 8'h44;
		memory[16'h18e8] <= 8'h6;
		memory[16'h18e9] <= 8'hb0;
		memory[16'h18ea] <= 8'h9d;
		memory[16'h18eb] <= 8'ha2;
		memory[16'h18ec] <= 8'h2;
		memory[16'h18ed] <= 8'haa;
		memory[16'h18ee] <= 8'h78;
		memory[16'h18ef] <= 8'haf;
		memory[16'h18f0] <= 8'ha1;
		memory[16'h18f1] <= 8'hcb;
		memory[16'h18f2] <= 8'hd6;
		memory[16'h18f3] <= 8'hcb;
		memory[16'h18f4] <= 8'he;
		memory[16'h18f5] <= 8'h7c;
		memory[16'h18f6] <= 8'h7b;
		memory[16'h18f7] <= 8'h83;
		memory[16'h18f8] <= 8'haa;
		memory[16'h18f9] <= 8'hc0;
		memory[16'h18fa] <= 8'h15;
		memory[16'h18fb] <= 8'h48;
		memory[16'h18fc] <= 8'hed;
		memory[16'h18fd] <= 8'h9f;
		memory[16'h18fe] <= 8'h5f;
		memory[16'h18ff] <= 8'h9c;
		memory[16'h1900] <= 8'h5b;
		memory[16'h1901] <= 8'h34;
		memory[16'h1902] <= 8'h36;
		memory[16'h1903] <= 8'h62;
		memory[16'h1904] <= 8'h38;
		memory[16'h1905] <= 8'h8e;
		memory[16'h1906] <= 8'ha7;
		memory[16'h1907] <= 8'h3e;
		memory[16'h1908] <= 8'h3e;
		memory[16'h1909] <= 8'h44;
		memory[16'h190a] <= 8'he0;
		memory[16'h190b] <= 8'h41;
		memory[16'h190c] <= 8'hee;
		memory[16'h190d] <= 8'h59;
		memory[16'h190e] <= 8'hf0;
		memory[16'h190f] <= 8'h8f;
		memory[16'h1910] <= 8'h24;
		memory[16'h1911] <= 8'hc6;
		memory[16'h1912] <= 8'h5b;
		memory[16'h1913] <= 8'h32;
		memory[16'h1914] <= 8'h43;
		memory[16'h1915] <= 8'hd6;
		memory[16'h1916] <= 8'hb5;
		memory[16'h1917] <= 8'hed;
		memory[16'h1918] <= 8'h96;
		memory[16'h1919] <= 8'hca;
		memory[16'h191a] <= 8'h35;
		memory[16'h191b] <= 8'h83;
		memory[16'h191c] <= 8'h6a;
		memory[16'h191d] <= 8'h95;
		memory[16'h191e] <= 8'h1f;
		memory[16'h191f] <= 8'hc5;
		memory[16'h1920] <= 8'hc9;
		memory[16'h1921] <= 8'h56;
		memory[16'h1922] <= 8'h28;
		memory[16'h1923] <= 8'h2;
		memory[16'h1924] <= 8'he4;
		memory[16'h1925] <= 8'hcf;
		memory[16'h1926] <= 8'h40;
		memory[16'h1927] <= 8'h23;
		memory[16'h1928] <= 8'h13;
		memory[16'h1929] <= 8'h21;
		memory[16'h192a] <= 8'h64;
		memory[16'h192b] <= 8'h1;
		memory[16'h192c] <= 8'h7a;
		memory[16'h192d] <= 8'h54;
		memory[16'h192e] <= 8'h90;
		memory[16'h192f] <= 8'h9e;
		memory[16'h1930] <= 8'h1a;
		memory[16'h1931] <= 8'heb;
		memory[16'h1932] <= 8'hd0;
		memory[16'h1933] <= 8'h5d;
		memory[16'h1934] <= 8'hc1;
		memory[16'h1935] <= 8'h85;
		memory[16'h1936] <= 8'h4a;
		memory[16'h1937] <= 8'h57;
		memory[16'h1938] <= 8'h50;
		memory[16'h1939] <= 8'h80;
		memory[16'h193a] <= 8'hda;
		memory[16'h193b] <= 8'hba;
		memory[16'h193c] <= 8'h15;
		memory[16'h193d] <= 8'hfa;
		memory[16'h193e] <= 8'h7f;
		memory[16'h193f] <= 8'hde;
		memory[16'h1940] <= 8'h50;
		memory[16'h1941] <= 8'ha7;
		memory[16'h1942] <= 8'he0;
		memory[16'h1943] <= 8'h34;
		memory[16'h1944] <= 8'h76;
		memory[16'h1945] <= 8'h21;
		memory[16'h1946] <= 8'h57;
		memory[16'h1947] <= 8'h89;
		memory[16'h1948] <= 8'h42;
		memory[16'h1949] <= 8'hbb;
		memory[16'h194a] <= 8'h8a;
		memory[16'h194b] <= 8'hbc;
		memory[16'h194c] <= 8'hf;
		memory[16'h194d] <= 8'h1b;
		memory[16'h194e] <= 8'h5a;
		memory[16'h194f] <= 8'h2a;
		memory[16'h1950] <= 8'h6;
		memory[16'h1951] <= 8'h2a;
		memory[16'h1952] <= 8'h87;
		memory[16'h1953] <= 8'hc8;
		memory[16'h1954] <= 8'haf;
		memory[16'h1955] <= 8'hd2;
		memory[16'h1956] <= 8'h1f;
		memory[16'h1957] <= 8'hff;
		memory[16'h1958] <= 8'h52;
		memory[16'h1959] <= 8'hfa;
		memory[16'h195a] <= 8'hb9;
		memory[16'h195b] <= 8'h67;
		memory[16'h195c] <= 8'hf4;
		memory[16'h195d] <= 8'h39;
		memory[16'h195e] <= 8'h45;
		memory[16'h195f] <= 8'h44;
		memory[16'h1960] <= 8'he0;
		memory[16'h1961] <= 8'h26;
		memory[16'h1962] <= 8'h78;
		memory[16'h1963] <= 8'h57;
		memory[16'h1964] <= 8'h47;
		memory[16'h1965] <= 8'hd0;
		memory[16'h1966] <= 8'he0;
		memory[16'h1967] <= 8'h89;
		memory[16'h1968] <= 8'h8b;
		memory[16'h1969] <= 8'h6b;
		memory[16'h196a] <= 8'h45;
		memory[16'h196b] <= 8'h9b;
		memory[16'h196c] <= 8'h86;
		memory[16'h196d] <= 8'h9f;
		memory[16'h196e] <= 8'hc5;
		memory[16'h196f] <= 8'h8c;
		memory[16'h1970] <= 8'hc9;
		memory[16'h1971] <= 8'h4c;
		memory[16'h1972] <= 8'h54;
		memory[16'h1973] <= 8'h78;
		memory[16'h1974] <= 8'h1e;
		memory[16'h1975] <= 8'h74;
		memory[16'h1976] <= 8'h78;
		memory[16'h1977] <= 8'h70;
		memory[16'h1978] <= 8'h6e;
		memory[16'h1979] <= 8'h31;
		memory[16'h197a] <= 8'hd7;
		memory[16'h197b] <= 8'h62;
		memory[16'h197c] <= 8'h6a;
		memory[16'h197d] <= 8'h1d;
		memory[16'h197e] <= 8'ha6;
		memory[16'h197f] <= 8'h4b;
		memory[16'h1980] <= 8'h43;
		memory[16'h1981] <= 8'h1e;
		memory[16'h1982] <= 8'ha2;
		memory[16'h1983] <= 8'h8a;
		memory[16'h1984] <= 8'hee;
		memory[16'h1985] <= 8'h82;
		memory[16'h1986] <= 8'h13;
		memory[16'h1987] <= 8'h7a;
		memory[16'h1988] <= 8'hed;
		memory[16'h1989] <= 8'h58;
		memory[16'h198a] <= 8'h15;
		memory[16'h198b] <= 8'h73;
		memory[16'h198c] <= 8'hf7;
		memory[16'h198d] <= 8'hda;
		memory[16'h198e] <= 8'h0;
		memory[16'h198f] <= 8'hc0;
		memory[16'h1990] <= 8'h26;
		memory[16'h1991] <= 8'h54;
		memory[16'h1992] <= 8'h38;
		memory[16'h1993] <= 8'h45;
		memory[16'h1994] <= 8'hc8;
		memory[16'h1995] <= 8'hb0;
		memory[16'h1996] <= 8'hb5;
		memory[16'h1997] <= 8'h36;
		memory[16'h1998] <= 8'he2;
		memory[16'h1999] <= 8'h8d;
		memory[16'h199a] <= 8'h98;
		memory[16'h199b] <= 8'h4c;
		memory[16'h199c] <= 8'haa;
		memory[16'h199d] <= 8'h3e;
		memory[16'h199e] <= 8'h97;
		memory[16'h199f] <= 8'hed;
		memory[16'h19a0] <= 8'h5d;
		memory[16'h19a1] <= 8'h39;
		memory[16'h19a2] <= 8'h77;
		memory[16'h19a3] <= 8'h4b;
		memory[16'h19a4] <= 8'hbc;
		memory[16'h19a5] <= 8'h8a;
		memory[16'h19a6] <= 8'hc5;
		memory[16'h19a7] <= 8'ha9;
		memory[16'h19a8] <= 8'he2;
		memory[16'h19a9] <= 8'hda;
		memory[16'h19aa] <= 8'h1d;
		memory[16'h19ab] <= 8'hd9;
		memory[16'h19ac] <= 8'hb4;
		memory[16'h19ad] <= 8'h1d;
		memory[16'h19ae] <= 8'h99;
		memory[16'h19af] <= 8'hdb;
		memory[16'h19b0] <= 8'h71;
		memory[16'h19b1] <= 8'hd1;
		memory[16'h19b2] <= 8'h20;
		memory[16'h19b3] <= 8'h3a;
		memory[16'h19b4] <= 8'h82;
		memory[16'h19b5] <= 8'hd5;
		memory[16'h19b6] <= 8'h70;
		memory[16'h19b7] <= 8'h64;
		memory[16'h19b8] <= 8'h62;
		memory[16'h19b9] <= 8'h9;
		memory[16'h19ba] <= 8'hb0;
		memory[16'h19bb] <= 8'hc;
		memory[16'h19bc] <= 8'h47;
		memory[16'h19bd] <= 8'h48;
		memory[16'h19be] <= 8'hf9;
		memory[16'h19bf] <= 8'ha4;
		memory[16'h19c0] <= 8'h81;
		memory[16'h19c1] <= 8'h70;
		memory[16'h19c2] <= 8'hf0;
		memory[16'h19c3] <= 8'h3d;
		memory[16'h19c4] <= 8'hfa;
		memory[16'h19c5] <= 8'hb5;
		memory[16'h19c6] <= 8'he7;
		memory[16'h19c7] <= 8'hdc;
		memory[16'h19c8] <= 8'h90;
		memory[16'h19c9] <= 8'h4;
		memory[16'h19ca] <= 8'hb5;
		memory[16'h19cb] <= 8'h44;
		memory[16'h19cc] <= 8'h21;
		memory[16'h19cd] <= 8'h4e;
		memory[16'h19ce] <= 8'h1f;
		memory[16'h19cf] <= 8'h92;
		memory[16'h19d0] <= 8'h20;
		memory[16'h19d1] <= 8'h3f;
		memory[16'h19d2] <= 8'hcc;
		memory[16'h19d3] <= 8'ha2;
		memory[16'h19d4] <= 8'h15;
		memory[16'h19d5] <= 8'h3d;
		memory[16'h19d6] <= 8'h6;
		memory[16'h19d7] <= 8'h77;
		memory[16'h19d8] <= 8'h46;
		memory[16'h19d9] <= 8'hb6;
		memory[16'h19da] <= 8'h84;
		memory[16'h19db] <= 8'h8d;
		memory[16'h19dc] <= 8'hfe;
		memory[16'h19dd] <= 8'h7d;
		memory[16'h19de] <= 8'h32;
		memory[16'h19df] <= 8'h80;
		memory[16'h19e0] <= 8'hee;
		memory[16'h19e1] <= 8'h22;
		memory[16'h19e2] <= 8'hbd;
		memory[16'h19e3] <= 8'he8;
		memory[16'h19e4] <= 8'hd7;
		memory[16'h19e5] <= 8'ha4;
		memory[16'h19e6] <= 8'hc5;
		memory[16'h19e7] <= 8'h67;
		memory[16'h19e8] <= 8'ha8;
		memory[16'h19e9] <= 8'h7a;
		memory[16'h19ea] <= 8'hac;
		memory[16'h19eb] <= 8'hc9;
		memory[16'h19ec] <= 8'hc9;
		memory[16'h19ed] <= 8'hcb;
		memory[16'h19ee] <= 8'h5c;
		memory[16'h19ef] <= 8'he9;
		memory[16'h19f0] <= 8'hb;
		memory[16'h19f1] <= 8'h28;
		memory[16'h19f2] <= 8'h8b;
		memory[16'h19f3] <= 8'h20;
		memory[16'h19f4] <= 8'h65;
		memory[16'h19f5] <= 8'h91;
		memory[16'h19f6] <= 8'h97;
		memory[16'h19f7] <= 8'hab;
		memory[16'h19f8] <= 8'h47;
		memory[16'h19f9] <= 8'h1b;
		memory[16'h19fa] <= 8'h39;
		memory[16'h19fb] <= 8'h46;
		memory[16'h19fc] <= 8'h99;
		memory[16'h19fd] <= 8'h6b;
		memory[16'h19fe] <= 8'hc6;
		memory[16'h19ff] <= 8'h87;
		memory[16'h1a00] <= 8'h8d;
		memory[16'h1a01] <= 8'h83;
		memory[16'h1a02] <= 8'h6f;
		memory[16'h1a03] <= 8'h64;
		memory[16'h1a04] <= 8'h28;
		memory[16'h1a05] <= 8'h34;
		memory[16'h1a06] <= 8'hcc;
		memory[16'h1a07] <= 8'hd0;
		memory[16'h1a08] <= 8'haf;
		memory[16'h1a09] <= 8'h78;
		memory[16'h1a0a] <= 8'h9a;
		memory[16'h1a0b] <= 8'h78;
		memory[16'h1a0c] <= 8'h43;
		memory[16'h1a0d] <= 8'hf6;
		memory[16'h1a0e] <= 8'h61;
		memory[16'h1a0f] <= 8'h4e;
		memory[16'h1a10] <= 8'h1e;
		memory[16'h1a11] <= 8'hec;
		memory[16'h1a12] <= 8'h6e;
		memory[16'h1a13] <= 8'h84;
		memory[16'h1a14] <= 8'h7d;
		memory[16'h1a15] <= 8'h6;
		memory[16'h1a16] <= 8'h2f;
		memory[16'h1a17] <= 8'hc4;
		memory[16'h1a18] <= 8'h21;
		memory[16'h1a19] <= 8'h68;
		memory[16'h1a1a] <= 8'ha;
		memory[16'h1a1b] <= 8'hba;
		memory[16'h1a1c] <= 8'hd3;
		memory[16'h1a1d] <= 8'hd0;
		memory[16'h1a1e] <= 8'h41;
		memory[16'h1a1f] <= 8'h60;
		memory[16'h1a20] <= 8'h54;
		memory[16'h1a21] <= 8'hb1;
		memory[16'h1a22] <= 8'hc5;
		memory[16'h1a23] <= 8'h7c;
		memory[16'h1a24] <= 8'he5;
		memory[16'h1a25] <= 8'h91;
		memory[16'h1a26] <= 8'h4c;
		memory[16'h1a27] <= 8'h94;
		memory[16'h1a28] <= 8'h9;
		memory[16'h1a29] <= 8'he6;
		memory[16'h1a2a] <= 8'hc;
		memory[16'h1a2b] <= 8'h4c;
		memory[16'h1a2c] <= 8'hdc;
		memory[16'h1a2d] <= 8'h6d;
		memory[16'h1a2e] <= 8'h9b;
		memory[16'h1a2f] <= 8'hfb;
		memory[16'h1a30] <= 8'h59;
		memory[16'h1a31] <= 8'h9;
		memory[16'h1a32] <= 8'h7f;
		memory[16'h1a33] <= 8'hd6;
		memory[16'h1a34] <= 8'hf;
		memory[16'h1a35] <= 8'hae;
		memory[16'h1a36] <= 8'h9b;
		memory[16'h1a37] <= 8'h31;
		memory[16'h1a38] <= 8'h17;
		memory[16'h1a39] <= 8'ha5;
		memory[16'h1a3a] <= 8'heb;
		memory[16'h1a3b] <= 8'hea;
		memory[16'h1a3c] <= 8'h76;
		memory[16'h1a3d] <= 8'h2d;
		memory[16'h1a3e] <= 8'h4b;
		memory[16'h1a3f] <= 8'hca;
		memory[16'h1a40] <= 8'hde;
		memory[16'h1a41] <= 8'h10;
		memory[16'h1a42] <= 8'h46;
		memory[16'h1a43] <= 8'hc3;
		memory[16'h1a44] <= 8'ha1;
		memory[16'h1a45] <= 8'h92;
		memory[16'h1a46] <= 8'h58;
		memory[16'h1a47] <= 8'haa;
		memory[16'h1a48] <= 8'h79;
		memory[16'h1a49] <= 8'h64;
		memory[16'h1a4a] <= 8'hf6;
		memory[16'h1a4b] <= 8'h55;
		memory[16'h1a4c] <= 8'hd2;
		memory[16'h1a4d] <= 8'h91;
		memory[16'h1a4e] <= 8'h50;
		memory[16'h1a4f] <= 8'h2b;
		memory[16'h1a50] <= 8'h9b;
		memory[16'h1a51] <= 8'hcf;
		memory[16'h1a52] <= 8'h2;
		memory[16'h1a53] <= 8'haa;
		memory[16'h1a54] <= 8'h7e;
		memory[16'h1a55] <= 8'h9d;
		memory[16'h1a56] <= 8'hdb;
		memory[16'h1a57] <= 8'h95;
		memory[16'h1a58] <= 8'h42;
		memory[16'h1a59] <= 8'hc7;
		memory[16'h1a5a] <= 8'h7f;
		memory[16'h1a5b] <= 8'hb8;
		memory[16'h1a5c] <= 8'hf4;
		memory[16'h1a5d] <= 8'hca;
		memory[16'h1a5e] <= 8'h82;
		memory[16'h1a5f] <= 8'hd2;
		memory[16'h1a60] <= 8'hda;
		memory[16'h1a61] <= 8'hc8;
		memory[16'h1a62] <= 8'h95;
		memory[16'h1a63] <= 8'h7b;
		memory[16'h1a64] <= 8'h5b;
		memory[16'h1a65] <= 8'hed;
		memory[16'h1a66] <= 8'h25;
		memory[16'h1a67] <= 8'hd4;
		memory[16'h1a68] <= 8'h52;
		memory[16'h1a69] <= 8'h1c;
		memory[16'h1a6a] <= 8'h29;
		memory[16'h1a6b] <= 8'h24;
		memory[16'h1a6c] <= 8'had;
		memory[16'h1a6d] <= 8'h7a;
		memory[16'h1a6e] <= 8'h4f;
		memory[16'h1a6f] <= 8'h48;
		memory[16'h1a70] <= 8'h49;
		memory[16'h1a71] <= 8'h51;
		memory[16'h1a72] <= 8'hf3;
		memory[16'h1a73] <= 8'hc7;
		memory[16'h1a74] <= 8'hee;
		memory[16'h1a75] <= 8'hce;
		memory[16'h1a76] <= 8'h5c;
		memory[16'h1a77] <= 8'h31;
		memory[16'h1a78] <= 8'h95;
		memory[16'h1a79] <= 8'hdc;
		memory[16'h1a7a] <= 8'he9;
		memory[16'h1a7b] <= 8'h89;
		memory[16'h1a7c] <= 8'ha6;
		memory[16'h1a7d] <= 8'h6c;
		memory[16'h1a7e] <= 8'h5b;
		memory[16'h1a7f] <= 8'h81;
		memory[16'h1a80] <= 8'h34;
		memory[16'h1a81] <= 8'hf1;
		memory[16'h1a82] <= 8'hfc;
		memory[16'h1a83] <= 8'h8f;
		memory[16'h1a84] <= 8'hde;
		memory[16'h1a85] <= 8'h22;
		memory[16'h1a86] <= 8'h63;
		memory[16'h1a87] <= 8'h30;
		memory[16'h1a88] <= 8'h3e;
		memory[16'h1a89] <= 8'h8d;
		memory[16'h1a8a] <= 8'h54;
		memory[16'h1a8b] <= 8'heb;
		memory[16'h1a8c] <= 8'h7;
		memory[16'h1a8d] <= 8'ha4;
		memory[16'h1a8e] <= 8'h34;
		memory[16'h1a8f] <= 8'h50;
		memory[16'h1a90] <= 8'hf5;
		memory[16'h1a91] <= 8'h27;
		memory[16'h1a92] <= 8'h18;
		memory[16'h1a93] <= 8'he4;
		memory[16'h1a94] <= 8'hf5;
		memory[16'h1a95] <= 8'h74;
		memory[16'h1a96] <= 8'h15;
		memory[16'h1a97] <= 8'h8b;
		memory[16'h1a98] <= 8'h50;
		memory[16'h1a99] <= 8'hfe;
		memory[16'h1a9a] <= 8'h14;
		memory[16'h1a9b] <= 8'hf7;
		memory[16'h1a9c] <= 8'h6a;
		memory[16'h1a9d] <= 8'h70;
		memory[16'h1a9e] <= 8'h78;
		memory[16'h1a9f] <= 8'h9f;
		memory[16'h1aa0] <= 8'h61;
		memory[16'h1aa1] <= 8'h74;
		memory[16'h1aa2] <= 8'h2e;
		memory[16'h1aa3] <= 8'h3f;
		memory[16'h1aa4] <= 8'h96;
		memory[16'h1aa5] <= 8'h92;
		memory[16'h1aa6] <= 8'h70;
		memory[16'h1aa7] <= 8'hd4;
		memory[16'h1aa8] <= 8'h1f;
		memory[16'h1aa9] <= 8'hc4;
		memory[16'h1aaa] <= 8'hc0;
		memory[16'h1aab] <= 8'h26;
		memory[16'h1aac] <= 8'h68;
		memory[16'h1aad] <= 8'hf4;
		memory[16'h1aae] <= 8'h76;
		memory[16'h1aaf] <= 8'h5e;
		memory[16'h1ab0] <= 8'h1b;
		memory[16'h1ab1] <= 8'h8e;
		memory[16'h1ab2] <= 8'h42;
		memory[16'h1ab3] <= 8'h10;
		memory[16'h1ab4] <= 8'h3;
		memory[16'h1ab5] <= 8'h57;
		memory[16'h1ab6] <= 8'h9b;
		memory[16'h1ab7] <= 8'h53;
		memory[16'h1ab8] <= 8'h55;
		memory[16'h1ab9] <= 8'hb0;
		memory[16'h1aba] <= 8'h4a;
		memory[16'h1abb] <= 8'hc0;
		memory[16'h1abc] <= 8'h20;
		memory[16'h1abd] <= 8'hc2;
		memory[16'h1abe] <= 8'h5f;
		memory[16'h1abf] <= 8'h81;
		memory[16'h1ac0] <= 8'h37;
		memory[16'h1ac1] <= 8'h8d;
		memory[16'h1ac2] <= 8'hc0;
		memory[16'h1ac3] <= 8'hcd;
		memory[16'h1ac4] <= 8'h1f;
		memory[16'h1ac5] <= 8'h30;
		memory[16'h1ac6] <= 8'ha2;
		memory[16'h1ac7] <= 8'h3e;
		memory[16'h1ac8] <= 8'hf5;
		memory[16'h1ac9] <= 8'h62;
		memory[16'h1aca] <= 8'h64;
		memory[16'h1acb] <= 8'h5d;
		memory[16'h1acc] <= 8'h56;
		memory[16'h1acd] <= 8'hdb;
		memory[16'h1ace] <= 8'hbb;
		memory[16'h1acf] <= 8'h71;
		memory[16'h1ad0] <= 8'h69;
		memory[16'h1ad1] <= 8'hfd;
		memory[16'h1ad2] <= 8'h81;
		memory[16'h1ad3] <= 8'h6c;
		memory[16'h1ad4] <= 8'h54;
		memory[16'h1ad5] <= 8'h1d;
		memory[16'h1ad6] <= 8'hc0;
		memory[16'h1ad7] <= 8'haa;
		memory[16'h1ad8] <= 8'hcd;
		memory[16'h1ad9] <= 8'ha;
		memory[16'h1ada] <= 8'h6a;
		memory[16'h1adb] <= 8'hed;
		memory[16'h1adc] <= 8'hcd;
		memory[16'h1add] <= 8'hc9;
		memory[16'h1ade] <= 8'h6e;
		memory[16'h1adf] <= 8'h4;
		memory[16'h1ae0] <= 8'h56;
		memory[16'h1ae1] <= 8'h2e;
		memory[16'h1ae2] <= 8'hd1;
		memory[16'h1ae3] <= 8'h76;
		memory[16'h1ae4] <= 8'h5f;
		memory[16'h1ae5] <= 8'h73;
		memory[16'h1ae6] <= 8'hb4;
		memory[16'h1ae7] <= 8'h54;
		memory[16'h1ae8] <= 8'hd5;
		memory[16'h1ae9] <= 8'h19;
		memory[16'h1aea] <= 8'hb1;
		memory[16'h1aeb] <= 8'h2b;
		memory[16'h1aec] <= 8'hf4;
		memory[16'h1aed] <= 8'h6d;
		memory[16'h1aee] <= 8'h9c;
		memory[16'h1aef] <= 8'h5d;
		memory[16'h1af0] <= 8'h6a;
		memory[16'h1af1] <= 8'h1e;
		memory[16'h1af2] <= 8'hca;
		memory[16'h1af3] <= 8'hbf;
		memory[16'h1af4] <= 8'h3b;
		memory[16'h1af5] <= 8'h8a;
		memory[16'h1af6] <= 8'h69;
		memory[16'h1af7] <= 8'h8;
		memory[16'h1af8] <= 8'h94;
		memory[16'h1af9] <= 8'hd3;
		memory[16'h1afa] <= 8'hf5;
		memory[16'h1afb] <= 8'h61;
		memory[16'h1afc] <= 8'h9c;
		memory[16'h1afd] <= 8'h63;
		memory[16'h1afe] <= 8'h65;
		memory[16'h1aff] <= 8'hf2;
		memory[16'h1b00] <= 8'h91;
		memory[16'h1b01] <= 8'h37;
		memory[16'h1b02] <= 8'h68;
		memory[16'h1b03] <= 8'hf0;
		memory[16'h1b04] <= 8'haa;
		memory[16'h1b05] <= 8'h1d;
		memory[16'h1b06] <= 8'h44;
		memory[16'h1b07] <= 8'h80;
		memory[16'h1b08] <= 8'h36;
		memory[16'h1b09] <= 8'hf6;
		memory[16'h1b0a] <= 8'hab;
		memory[16'h1b0b] <= 8'h2a;
		memory[16'h1b0c] <= 8'h63;
		memory[16'h1b0d] <= 8'h48;
		memory[16'h1b0e] <= 8'h87;
		memory[16'h1b0f] <= 8'hcd;
		memory[16'h1b10] <= 8'h66;
		memory[16'h1b11] <= 8'h51;
		memory[16'h1b12] <= 8'h8c;
		memory[16'h1b13] <= 8'ha1;
		memory[16'h1b14] <= 8'hdb;
		memory[16'h1b15] <= 8'hf5;
		memory[16'h1b16] <= 8'ha9;
		memory[16'h1b17] <= 8'h70;
		memory[16'h1b18] <= 8'hc8;
		memory[16'h1b19] <= 8'h9e;
		memory[16'h1b1a] <= 8'hd1;
		memory[16'h1b1b] <= 8'h64;
		memory[16'h1b1c] <= 8'h1;
		memory[16'h1b1d] <= 8'h37;
		memory[16'h1b1e] <= 8'h57;
		memory[16'h1b1f] <= 8'h92;
		memory[16'h1b20] <= 8'h6e;
		memory[16'h1b21] <= 8'hbf;
		memory[16'h1b22] <= 8'h83;
		memory[16'h1b23] <= 8'h18;
		memory[16'h1b24] <= 8'hdc;
		memory[16'h1b25] <= 8'hc7;
		memory[16'h1b26] <= 8'h98;
		memory[16'h1b27] <= 8'h12;
		memory[16'h1b28] <= 8'hbd;
		memory[16'h1b29] <= 8'h44;
		memory[16'h1b2a] <= 8'h3c;
		memory[16'h1b2b] <= 8'h20;
		memory[16'h1b2c] <= 8'h8c;
		memory[16'h1b2d] <= 8'hc4;
		memory[16'h1b2e] <= 8'hee;
		memory[16'h1b2f] <= 8'hf2;
		memory[16'h1b30] <= 8'h15;
		memory[16'h1b31] <= 8'h7a;
		memory[16'h1b32] <= 8'h93;
		memory[16'h1b33] <= 8'hf1;
		memory[16'h1b34] <= 8'h70;
		memory[16'h1b35] <= 8'h3c;
		memory[16'h1b36] <= 8'h61;
		memory[16'h1b37] <= 8'h38;
		memory[16'h1b38] <= 8'hda;
		memory[16'h1b39] <= 8'h32;
		memory[16'h1b3a] <= 8'h9d;
		memory[16'h1b3b] <= 8'hdb;
		memory[16'h1b3c] <= 8'h69;
		memory[16'h1b3d] <= 8'hf4;
		memory[16'h1b3e] <= 8'h6d;
		memory[16'h1b3f] <= 8'hd7;
		memory[16'h1b40] <= 8'hb3;
		memory[16'h1b41] <= 8'hf0;
		memory[16'h1b42] <= 8'hf0;
		memory[16'h1b43] <= 8'h90;
		memory[16'h1b44] <= 8'hb8;
		memory[16'h1b45] <= 8'h88;
		memory[16'h1b46] <= 8'ha2;
		memory[16'h1b47] <= 8'h75;
		memory[16'h1b48] <= 8'hcc;
		memory[16'h1b49] <= 8'hdf;
		memory[16'h1b4a] <= 8'h96;
		memory[16'h1b4b] <= 8'h58;
		memory[16'h1b4c] <= 8'ha3;
		memory[16'h1b4d] <= 8'h84;
		memory[16'h1b4e] <= 8'h4a;
		memory[16'h1b4f] <= 8'hb8;
		memory[16'h1b50] <= 8'hfe;
		memory[16'h1b51] <= 8'hdd;
		memory[16'h1b52] <= 8'ha9;
		memory[16'h1b53] <= 8'h6e;
		memory[16'h1b54] <= 8'h19;
		memory[16'h1b55] <= 8'ha;
		memory[16'h1b56] <= 8'ha7;
		memory[16'h1b57] <= 8'hf3;
		memory[16'h1b58] <= 8'h3d;
		memory[16'h1b59] <= 8'h44;
		memory[16'h1b5a] <= 8'hce;
		memory[16'h1b5b] <= 8'ha6;
		memory[16'h1b5c] <= 8'h38;
		memory[16'h1b5d] <= 8'h3c;
		memory[16'h1b5e] <= 8'h7e;
		memory[16'h1b5f] <= 8'heb;
		memory[16'h1b60] <= 8'h2c;
		memory[16'h1b61] <= 8'h6e;
		memory[16'h1b62] <= 8'h7b;
		memory[16'h1b63] <= 8'he4;
		memory[16'h1b64] <= 8'hf6;
		memory[16'h1b65] <= 8'h1e;
		memory[16'h1b66] <= 8'h5a;
		memory[16'h1b67] <= 8'hc3;
		memory[16'h1b68] <= 8'hfd;
		memory[16'h1b69] <= 8'hf0;
		memory[16'h1b6a] <= 8'h1b;
		memory[16'h1b6b] <= 8'ha0;
		memory[16'h1b6c] <= 8'h74;
		memory[16'h1b6d] <= 8'h66;
		memory[16'h1b6e] <= 8'h58;
		memory[16'h1b6f] <= 8'h72;
		memory[16'h1b70] <= 8'h43;
		memory[16'h1b71] <= 8'h2;
		memory[16'h1b72] <= 8'he1;
		memory[16'h1b73] <= 8'h5d;
		memory[16'h1b74] <= 8'hc;
		memory[16'h1b75] <= 8'h88;
		memory[16'h1b76] <= 8'h50;
		memory[16'h1b77] <= 8'h49;
		memory[16'h1b78] <= 8'hcc;
		memory[16'h1b79] <= 8'h1f;
		memory[16'h1b7a] <= 8'hf0;
		memory[16'h1b7b] <= 8'h4;
		memory[16'h1b7c] <= 8'h5b;
		memory[16'h1b7d] <= 8'h6e;
		memory[16'h1b7e] <= 8'hef;
		memory[16'h1b7f] <= 8'h87;
		memory[16'h1b80] <= 8'hdc;
		memory[16'h1b81] <= 8'h6b;
		memory[16'h1b82] <= 8'h6c;
		memory[16'h1b83] <= 8'hd2;
		memory[16'h1b84] <= 8'h89;
		memory[16'h1b85] <= 8'hc6;
		memory[16'h1b86] <= 8'h95;
		memory[16'h1b87] <= 8'h86;
		memory[16'h1b88] <= 8'hb6;
		memory[16'h1b89] <= 8'hb1;
		memory[16'h1b8a] <= 8'h26;
		memory[16'h1b8b] <= 8'h2a;
		memory[16'h1b8c] <= 8'h17;
		memory[16'h1b8d] <= 8'h7e;
		memory[16'h1b8e] <= 8'h9c;
		memory[16'h1b8f] <= 8'h5a;
		memory[16'h1b90] <= 8'h80;
		memory[16'h1b91] <= 8'h7d;
		memory[16'h1b92] <= 8'hb7;
		memory[16'h1b93] <= 8'h8d;
		memory[16'h1b94] <= 8'h5;
		memory[16'h1b95] <= 8'h8;
		memory[16'h1b96] <= 8'hd6;
		memory[16'h1b97] <= 8'hd1;
		memory[16'h1b98] <= 8'h27;
		memory[16'h1b99] <= 8'hc6;
		memory[16'h1b9a] <= 8'hd5;
		memory[16'h1b9b] <= 8'h82;
		memory[16'h1b9c] <= 8'h34;
		memory[16'h1b9d] <= 8'hc5;
		memory[16'h1b9e] <= 8'h9;
		memory[16'h1b9f] <= 8'h10;
		memory[16'h1ba0] <= 8'h30;
		memory[16'h1ba1] <= 8'h75;
		memory[16'h1ba2] <= 8'he3;
		memory[16'h1ba3] <= 8'hb9;
		memory[16'h1ba4] <= 8'h3b;
		memory[16'h1ba5] <= 8'h78;
		memory[16'h1ba6] <= 8'h3f;
		memory[16'h1ba7] <= 8'hf1;
		memory[16'h1ba8] <= 8'h29;
		memory[16'h1ba9] <= 8'h65;
		memory[16'h1baa] <= 8'h1b;
		memory[16'h1bab] <= 8'h40;
		memory[16'h1bac] <= 8'he3;
		memory[16'h1bad] <= 8'hb8;
		memory[16'h1bae] <= 8'h9b;
		memory[16'h1baf] <= 8'h64;
		memory[16'h1bb0] <= 8'h35;
		memory[16'h1bb1] <= 8'h52;
		memory[16'h1bb2] <= 8'hf1;
		memory[16'h1bb3] <= 8'h3b;
		memory[16'h1bb4] <= 8'h5a;
		memory[16'h1bb5] <= 8'hc7;
		memory[16'h1bb6] <= 8'hc;
		memory[16'h1bb7] <= 8'h81;
		memory[16'h1bb8] <= 8'h8e;
		memory[16'h1bb9] <= 8'he2;
		memory[16'h1bba] <= 8'h3;
		memory[16'h1bbb] <= 8'hc2;
		memory[16'h1bbc] <= 8'ha7;
		memory[16'h1bbd] <= 8'hd;
		memory[16'h1bbe] <= 8'hd3;
		memory[16'h1bbf] <= 8'hd7;
		memory[16'h1bc0] <= 8'h82;
		memory[16'h1bc1] <= 8'hb6;
		memory[16'h1bc2] <= 8'h90;
		memory[16'h1bc3] <= 8'hbe;
		memory[16'h1bc4] <= 8'h2e;
		memory[16'h1bc5] <= 8'hcf;
		memory[16'h1bc6] <= 8'haf;
		memory[16'h1bc7] <= 8'h58;
		memory[16'h1bc8] <= 8'h34;
		memory[16'h1bc9] <= 8'hcb;
		memory[16'h1bca] <= 8'h98;
		memory[16'h1bcb] <= 8'h17;
		memory[16'h1bcc] <= 8'h83;
		memory[16'h1bcd] <= 8'h33;
		memory[16'h1bce] <= 8'h7b;
		memory[16'h1bcf] <= 8'hb8;
		memory[16'h1bd0] <= 8'h86;
		memory[16'h1bd1] <= 8'h6c;
		memory[16'h1bd2] <= 8'hf3;
		memory[16'h1bd3] <= 8'he0;
		memory[16'h1bd4] <= 8'h34;
		memory[16'h1bd5] <= 8'h0;
		memory[16'h1bd6] <= 8'h62;
		memory[16'h1bd7] <= 8'hc2;
		memory[16'h1bd8] <= 8'he2;
		memory[16'h1bd9] <= 8'h65;
		memory[16'h1bda] <= 8'h84;
		memory[16'h1bdb] <= 8'h89;
		memory[16'h1bdc] <= 8'h72;
		memory[16'h1bdd] <= 8'h57;
		memory[16'h1bde] <= 8'h60;
		memory[16'h1bdf] <= 8'hf5;
		memory[16'h1be0] <= 8'hd;
		memory[16'h1be1] <= 8'hf0;
		memory[16'h1be2] <= 8'hb3;
		memory[16'h1be3] <= 8'h3c;
		memory[16'h1be4] <= 8'hbf;
		memory[16'h1be5] <= 8'h62;
		memory[16'h1be6] <= 8'h94;
		memory[16'h1be7] <= 8'hf3;
		memory[16'h1be8] <= 8'h2d;
		memory[16'h1be9] <= 8'h2c;
		memory[16'h1bea] <= 8'ha;
		memory[16'h1beb] <= 8'hb0;
		memory[16'h1bec] <= 8'h60;
		memory[16'h1bed] <= 8'h86;
		memory[16'h1bee] <= 8'h69;
		memory[16'h1bef] <= 8'he6;
		memory[16'h1bf0] <= 8'hf2;
		memory[16'h1bf1] <= 8'h5c;
		memory[16'h1bf2] <= 8'hc6;
		memory[16'h1bf3] <= 8'h26;
		memory[16'h1bf4] <= 8'h5c;
		memory[16'h1bf5] <= 8'h28;
		memory[16'h1bf6] <= 8'he8;
		memory[16'h1bf7] <= 8'h3e;
		memory[16'h1bf8] <= 8'h8e;
		memory[16'h1bf9] <= 8'h6d;
		memory[16'h1bfa] <= 8'hc7;
		memory[16'h1bfb] <= 8'h0;
		memory[16'h1bfc] <= 8'hc4;
		memory[16'h1bfd] <= 8'h27;
		memory[16'h1bfe] <= 8'hf5;
		memory[16'h1bff] <= 8'hd2;
		memory[16'h1c00] <= 8'h17;
		memory[16'h1c01] <= 8'ha8;
		memory[16'h1c02] <= 8'he;
		memory[16'h1c03] <= 8'hd6;
		memory[16'h1c04] <= 8'hb;
		memory[16'h1c05] <= 8'ha2;
		memory[16'h1c06] <= 8'hc9;
		memory[16'h1c07] <= 8'h38;
		memory[16'h1c08] <= 8'hce;
		memory[16'h1c09] <= 8'hd4;
		memory[16'h1c0a] <= 8'he9;
		memory[16'h1c0b] <= 8'h2e;
		memory[16'h1c0c] <= 8'h5a;
		memory[16'h1c0d] <= 8'h52;
		memory[16'h1c0e] <= 8'h14;
		memory[16'h1c0f] <= 8'h4c;
		memory[16'h1c10] <= 8'hae;
		memory[16'h1c11] <= 8'hdb;
		memory[16'h1c12] <= 8'h73;
		memory[16'h1c13] <= 8'hb;
		memory[16'h1c14] <= 8'h3;
		memory[16'h1c15] <= 8'h5b;
		memory[16'h1c16] <= 8'h49;
		memory[16'h1c17] <= 8'h91;
		memory[16'h1c18] <= 8'hc8;
		memory[16'h1c19] <= 8'h11;
		memory[16'h1c1a] <= 8'h92;
		memory[16'h1c1b] <= 8'h8d;
		memory[16'h1c1c] <= 8'h38;
		memory[16'h1c1d] <= 8'h87;
		memory[16'h1c1e] <= 8'h5f;
		memory[16'h1c1f] <= 8'h50;
		memory[16'h1c20] <= 8'h30;
		memory[16'h1c21] <= 8'h6d;
		memory[16'h1c22] <= 8'h26;
		memory[16'h1c23] <= 8'h3b;
		memory[16'h1c24] <= 8'hf;
		memory[16'h1c25] <= 8'hf0;
		memory[16'h1c26] <= 8'h73;
		memory[16'h1c27] <= 8'hdd;
		memory[16'h1c28] <= 8'hc4;
		memory[16'h1c29] <= 8'h5c;
		memory[16'h1c2a] <= 8'hc;
		memory[16'h1c2b] <= 8'h1e;
		memory[16'h1c2c] <= 8'hae;
		memory[16'h1c2d] <= 8'h20;
		memory[16'h1c2e] <= 8'h6a;
		memory[16'h1c2f] <= 8'h5d;
		memory[16'h1c30] <= 8'hfb;
		memory[16'h1c31] <= 8'hdd;
		memory[16'h1c32] <= 8'h68;
		memory[16'h1c33] <= 8'hff;
		memory[16'h1c34] <= 8'h39;
		memory[16'h1c35] <= 8'hb1;
		memory[16'h1c36] <= 8'h90;
		memory[16'h1c37] <= 8'h1;
		memory[16'h1c38] <= 8'hc2;
		memory[16'h1c39] <= 8'h22;
		memory[16'h1c3a] <= 8'h8e;
		memory[16'h1c3b] <= 8'hfb;
		memory[16'h1c3c] <= 8'haa;
		memory[16'h1c3d] <= 8'hed;
		memory[16'h1c3e] <= 8'h4b;
		memory[16'h1c3f] <= 8'hda;
		memory[16'h1c40] <= 8'h5a;
		memory[16'h1c41] <= 8'h71;
		memory[16'h1c42] <= 8'h15;
		memory[16'h1c43] <= 8'h69;
		memory[16'h1c44] <= 8'h61;
		memory[16'h1c45] <= 8'h88;
		memory[16'h1c46] <= 8'h47;
		memory[16'h1c47] <= 8'h25;
		memory[16'h1c48] <= 8'he5;
		memory[16'h1c49] <= 8'h53;
		memory[16'h1c4a] <= 8'h43;
		memory[16'h1c4b] <= 8'h93;
		memory[16'h1c4c] <= 8'h73;
		memory[16'h1c4d] <= 8'hae;
		memory[16'h1c4e] <= 8'hf0;
		memory[16'h1c4f] <= 8'h6f;
		memory[16'h1c50] <= 8'h8b;
		memory[16'h1c51] <= 8'h58;
		memory[16'h1c52] <= 8'h6e;
		memory[16'h1c53] <= 8'hc4;
		memory[16'h1c54] <= 8'ha;
		memory[16'h1c55] <= 8'hfe;
		memory[16'h1c56] <= 8'hc6;
		memory[16'h1c57] <= 8'hcc;
		memory[16'h1c58] <= 8'h21;
		memory[16'h1c59] <= 8'h54;
		memory[16'h1c5a] <= 8'hc7;
		memory[16'h1c5b] <= 8'hcb;
		memory[16'h1c5c] <= 8'h42;
		memory[16'h1c5d] <= 8'h12;
		memory[16'h1c5e] <= 8'ha5;
		memory[16'h1c5f] <= 8'h9c;
		memory[16'h1c60] <= 8'h84;
		memory[16'h1c61] <= 8'hba;
		memory[16'h1c62] <= 8'h6;
		memory[16'h1c63] <= 8'he5;
		memory[16'h1c64] <= 8'h42;
		memory[16'h1c65] <= 8'h4d;
		memory[16'h1c66] <= 8'hb;
		memory[16'h1c67] <= 8'h27;
		memory[16'h1c68] <= 8'ha0;
		memory[16'h1c69] <= 8'h4e;
		memory[16'h1c6a] <= 8'hbb;
		memory[16'h1c6b] <= 8'h13;
		memory[16'h1c6c] <= 8'hfc;
		memory[16'h1c6d] <= 8'hab;
		memory[16'h1c6e] <= 8'h82;
		memory[16'h1c6f] <= 8'h88;
		memory[16'h1c70] <= 8'h4;
		memory[16'h1c71] <= 8'hf0;
		memory[16'h1c72] <= 8'h4c;
		memory[16'h1c73] <= 8'he;
		memory[16'h1c74] <= 8'hef;
		memory[16'h1c75] <= 8'h12;
		memory[16'h1c76] <= 8'hda;
		memory[16'h1c77] <= 8'h10;
		memory[16'h1c78] <= 8'h67;
		memory[16'h1c79] <= 8'ha2;
		memory[16'h1c7a] <= 8'hdb;
		memory[16'h1c7b] <= 8'ha9;
		memory[16'h1c7c] <= 8'hb4;
		memory[16'h1c7d] <= 8'h80;
		memory[16'h1c7e] <= 8'h45;
		memory[16'h1c7f] <= 8'h38;
		memory[16'h1c80] <= 8'h3a;
		memory[16'h1c81] <= 8'h4b;
		memory[16'h1c82] <= 8'h1e;
		memory[16'h1c83] <= 8'h7c;
		memory[16'h1c84] <= 8'h98;
		memory[16'h1c85] <= 8'h29;
		memory[16'h1c86] <= 8'ha4;
		memory[16'h1c87] <= 8'h38;
		memory[16'h1c88] <= 8'h77;
		memory[16'h1c89] <= 8'h5f;
		memory[16'h1c8a] <= 8'h4c;
		memory[16'h1c8b] <= 8'h74;
		memory[16'h1c8c] <= 8'ha;
		memory[16'h1c8d] <= 8'hce;
		memory[16'h1c8e] <= 8'hfc;
		memory[16'h1c8f] <= 8'he;
		memory[16'h1c90] <= 8'hbf;
		memory[16'h1c91] <= 8'h48;
		memory[16'h1c92] <= 8'h1c;
		memory[16'h1c93] <= 8'hae;
		memory[16'h1c94] <= 8'h5b;
		memory[16'h1c95] <= 8'hf7;
		memory[16'h1c96] <= 8'hbe;
		memory[16'h1c97] <= 8'hc2;
		memory[16'h1c98] <= 8'h99;
		memory[16'h1c99] <= 8'h99;
		memory[16'h1c9a] <= 8'h6b;
		memory[16'h1c9b] <= 8'h4d;
		memory[16'h1c9c] <= 8'h19;
		memory[16'h1c9d] <= 8'hb0;
		memory[16'h1c9e] <= 8'h86;
		memory[16'h1c9f] <= 8'h53;
		memory[16'h1ca0] <= 8'hfc;
		memory[16'h1ca1] <= 8'ha4;
		memory[16'h1ca2] <= 8'hcf;
		memory[16'h1ca3] <= 8'h94;
		memory[16'h1ca4] <= 8'hcd;
		memory[16'h1ca5] <= 8'h73;
		memory[16'h1ca6] <= 8'hcd;
		memory[16'h1ca7] <= 8'h44;
		memory[16'h1ca8] <= 8'hd2;
		memory[16'h1ca9] <= 8'h19;
		memory[16'h1caa] <= 8'hb8;
		memory[16'h1cab] <= 8'hdd;
		memory[16'h1cac] <= 8'he7;
		memory[16'h1cad] <= 8'hb4;
		memory[16'h1cae] <= 8'heb;
		memory[16'h1caf] <= 8'ha6;
		memory[16'h1cb0] <= 8'hfd;
		memory[16'h1cb1] <= 8'h8;
		memory[16'h1cb2] <= 8'h54;
		memory[16'h1cb3] <= 8'h58;
		memory[16'h1cb4] <= 8'hff;
		memory[16'h1cb5] <= 8'h12;
		memory[16'h1cb6] <= 8'h1a;
		memory[16'h1cb7] <= 8'h98;
		memory[16'h1cb8] <= 8'hab;
		memory[16'h1cb9] <= 8'h85;
		memory[16'h1cba] <= 8'he5;
		memory[16'h1cbb] <= 8'hc4;
		memory[16'h1cbc] <= 8'h35;
		memory[16'h1cbd] <= 8'h6b;
		memory[16'h1cbe] <= 8'h17;
		memory[16'h1cbf] <= 8'h31;
		memory[16'h1cc0] <= 8'hf;
		memory[16'h1cc1] <= 8'he7;
		memory[16'h1cc2] <= 8'hc6;
		memory[16'h1cc3] <= 8'hdc;
		memory[16'h1cc4] <= 8'h5a;
		memory[16'h1cc5] <= 8'h93;
		memory[16'h1cc6] <= 8'h21;
		memory[16'h1cc7] <= 8'h2d;
		memory[16'h1cc8] <= 8'hac;
		memory[16'h1cc9] <= 8'hd9;
		memory[16'h1cca] <= 8'ha;
		memory[16'h1ccb] <= 8'h93;
		memory[16'h1ccc] <= 8'h8e;
		memory[16'h1ccd] <= 8'hf5;
		memory[16'h1cce] <= 8'h3a;
		memory[16'h1ccf] <= 8'h8b;
		memory[16'h1cd0] <= 8'hfd;
		memory[16'h1cd1] <= 8'h8e;
		memory[16'h1cd2] <= 8'he3;
		memory[16'h1cd3] <= 8'hfc;
		memory[16'h1cd4] <= 8'ha1;
		memory[16'h1cd5] <= 8'hfd;
		memory[16'h1cd6] <= 8'h94;
		memory[16'h1cd7] <= 8'h4c;
		memory[16'h1cd8] <= 8'h82;
		memory[16'h1cd9] <= 8'h7a;
		memory[16'h1cda] <= 8'h11;
		memory[16'h1cdb] <= 8'hb7;
		memory[16'h1cdc] <= 8'he5;
		memory[16'h1cdd] <= 8'h28;
		memory[16'h1cde] <= 8'he9;
		memory[16'h1cdf] <= 8'hf5;
		memory[16'h1ce0] <= 8'hf;
		memory[16'h1ce1] <= 8'haf;
		memory[16'h1ce2] <= 8'hd1;
		memory[16'h1ce3] <= 8'h6a;
		memory[16'h1ce4] <= 8'h42;
		memory[16'h1ce5] <= 8'hf2;
		memory[16'h1ce6] <= 8'h97;
		memory[16'h1ce7] <= 8'hee;
		memory[16'h1ce8] <= 8'hcc;
		memory[16'h1ce9] <= 8'ha1;
		memory[16'h1cea] <= 8'h81;
		memory[16'h1ceb] <= 8'h5a;
		memory[16'h1cec] <= 8'h96;
		memory[16'h1ced] <= 8'hbb;
		memory[16'h1cee] <= 8'he5;
		memory[16'h1cef] <= 8'h94;
		memory[16'h1cf0] <= 8'h4a;
		memory[16'h1cf1] <= 8'hc8;
		memory[16'h1cf2] <= 8'h90;
		memory[16'h1cf3] <= 8'heb;
		memory[16'h1cf4] <= 8'hc5;
		memory[16'h1cf5] <= 8'h25;
		memory[16'h1cf6] <= 8'h37;
		memory[16'h1cf7] <= 8'h47;
		memory[16'h1cf8] <= 8'h9f;
		memory[16'h1cf9] <= 8'h48;
		memory[16'h1cfa] <= 8'hfe;
		memory[16'h1cfb] <= 8'h84;
		memory[16'h1cfc] <= 8'h71;
		memory[16'h1cfd] <= 8'he7;
		memory[16'h1cfe] <= 8'h79;
		memory[16'h1cff] <= 8'h80;
		memory[16'h1d00] <= 8'h96;
		memory[16'h1d01] <= 8'h4b;
		memory[16'h1d02] <= 8'hea;
		memory[16'h1d03] <= 8'hd8;
		memory[16'h1d04] <= 8'h3d;
		memory[16'h1d05] <= 8'h81;
		memory[16'h1d06] <= 8'hc6;
		memory[16'h1d07] <= 8'h9;
		memory[16'h1d08] <= 8'h22;
		memory[16'h1d09] <= 8'h48;
		memory[16'h1d0a] <= 8'h63;
		memory[16'h1d0b] <= 8'hb9;
		memory[16'h1d0c] <= 8'h3;
		memory[16'h1d0d] <= 8'h48;
		memory[16'h1d0e] <= 8'h4d;
		memory[16'h1d0f] <= 8'h4d;
		memory[16'h1d10] <= 8'h10;
		memory[16'h1d11] <= 8'hdd;
		memory[16'h1d12] <= 8'h38;
		memory[16'h1d13] <= 8'hd5;
		memory[16'h1d14] <= 8'h2;
		memory[16'h1d15] <= 8'h70;
		memory[16'h1d16] <= 8'h1c;
		memory[16'h1d17] <= 8'ha1;
		memory[16'h1d18] <= 8'hb8;
		memory[16'h1d19] <= 8'h1b;
		memory[16'h1d1a] <= 8'h26;
		memory[16'h1d1b] <= 8'h29;
		memory[16'h1d1c] <= 8'h2;
		memory[16'h1d1d] <= 8'h9f;
		memory[16'h1d1e] <= 8'haa;
		memory[16'h1d1f] <= 8'h99;
		memory[16'h1d20] <= 8'hea;
		memory[16'h1d21] <= 8'h94;
		memory[16'h1d22] <= 8'h71;
		memory[16'h1d23] <= 8'h28;
		memory[16'h1d24] <= 8'h16;
		memory[16'h1d25] <= 8'h38;
		memory[16'h1d26] <= 8'h31;
		memory[16'h1d27] <= 8'h38;
		memory[16'h1d28] <= 8'h80;
		memory[16'h1d29] <= 8'h95;
		memory[16'h1d2a] <= 8'hf1;
		memory[16'h1d2b] <= 8'h83;
		memory[16'h1d2c] <= 8'hdd;
		memory[16'h1d2d] <= 8'h3e;
		memory[16'h1d2e] <= 8'hd1;
		memory[16'h1d2f] <= 8'hee;
		memory[16'h1d30] <= 8'h1c;
		memory[16'h1d31] <= 8'h9;
		memory[16'h1d32] <= 8'hc3;
		memory[16'h1d33] <= 8'h1e;
		memory[16'h1d34] <= 8'h79;
		memory[16'h1d35] <= 8'he0;
		memory[16'h1d36] <= 8'hc0;
		memory[16'h1d37] <= 8'h32;
		memory[16'h1d38] <= 8'hfb;
		memory[16'h1d39] <= 8'he6;
		memory[16'h1d3a] <= 8'h5b;
		memory[16'h1d3b] <= 8'hfd;
		memory[16'h1d3c] <= 8'h85;
		memory[16'h1d3d] <= 8'h5;
		memory[16'h1d3e] <= 8'h96;
		memory[16'h1d3f] <= 8'h70;
		memory[16'h1d40] <= 8'h9a;
		memory[16'h1d41] <= 8'h8;
		memory[16'h1d42] <= 8'h98;
		memory[16'h1d43] <= 8'hb0;
		memory[16'h1d44] <= 8'h40;
		memory[16'h1d45] <= 8'hc9;
		memory[16'h1d46] <= 8'he8;
		memory[16'h1d47] <= 8'hc0;
		memory[16'h1d48] <= 8'h5e;
		memory[16'h1d49] <= 8'hda;
		memory[16'h1d4a] <= 8'h43;
		memory[16'h1d4b] <= 8'h3c;
		memory[16'h1d4c] <= 8'h18;
		memory[16'h1d4d] <= 8'h14;
		memory[16'h1d4e] <= 8'h2a;
		memory[16'h1d4f] <= 8'h34;
		memory[16'h1d50] <= 8'h1e;
		memory[16'h1d51] <= 8'hed;
		memory[16'h1d52] <= 8'h53;
		memory[16'h1d53] <= 8'h97;
		memory[16'h1d54] <= 8'hcd;
		memory[16'h1d55] <= 8'h13;
		memory[16'h1d56] <= 8'hc9;
		memory[16'h1d57] <= 8'hc8;
		memory[16'h1d58] <= 8'hf9;
		memory[16'h1d59] <= 8'h25;
		memory[16'h1d5a] <= 8'hc6;
		memory[16'h1d5b] <= 8'h7e;
		memory[16'h1d5c] <= 8'h2a;
		memory[16'h1d5d] <= 8'h5c;
		memory[16'h1d5e] <= 8'hee;
		memory[16'h1d5f] <= 8'hc4;
		memory[16'h1d60] <= 8'h64;
		memory[16'h1d61] <= 8'h86;
		memory[16'h1d62] <= 8'h74;
		memory[16'h1d63] <= 8'ha4;
		memory[16'h1d64] <= 8'h50;
		memory[16'h1d65] <= 8'h5d;
		memory[16'h1d66] <= 8'h64;
		memory[16'h1d67] <= 8'hae;
		memory[16'h1d68] <= 8'h37;
		memory[16'h1d69] <= 8'ha8;
		memory[16'h1d6a] <= 8'hea;
		memory[16'h1d6b] <= 8'h4f;
		memory[16'h1d6c] <= 8'hbc;
		memory[16'h1d6d] <= 8'h14;
		memory[16'h1d6e] <= 8'h84;
		memory[16'h1d6f] <= 8'hda;
		memory[16'h1d70] <= 8'h2;
		memory[16'h1d71] <= 8'hd7;
		memory[16'h1d72] <= 8'h72;
		memory[16'h1d73] <= 8'hcf;
		memory[16'h1d74] <= 8'hea;
		memory[16'h1d75] <= 8'h3b;
		memory[16'h1d76] <= 8'h98;
		memory[16'h1d77] <= 8'he3;
		memory[16'h1d78] <= 8'h60;
		memory[16'h1d79] <= 8'h5e;
		memory[16'h1d7a] <= 8'h61;
		memory[16'h1d7b] <= 8'h8b;
		memory[16'h1d7c] <= 8'hba;
		memory[16'h1d7d] <= 8'h50;
		memory[16'h1d7e] <= 8'h4f;
		memory[16'h1d7f] <= 8'h1f;
		memory[16'h1d80] <= 8'hd6;
		memory[16'h1d81] <= 8'hc4;
		memory[16'h1d82] <= 8'hc3;
		memory[16'h1d83] <= 8'h26;
		memory[16'h1d84] <= 8'h21;
		memory[16'h1d85] <= 8'h28;
		memory[16'h1d86] <= 8'hd5;
		memory[16'h1d87] <= 8'h58;
		memory[16'h1d88] <= 8'hd0;
		memory[16'h1d89] <= 8'hbf;
		memory[16'h1d8a] <= 8'ha7;
		memory[16'h1d8b] <= 8'h8c;
		memory[16'h1d8c] <= 8'hd4;
		memory[16'h1d8d] <= 8'h2b;
		memory[16'h1d8e] <= 8'h67;
		memory[16'h1d8f] <= 8'hd6;
		memory[16'h1d90] <= 8'h2;
		memory[16'h1d91] <= 8'hd9;
		memory[16'h1d92] <= 8'ha5;
		memory[16'h1d93] <= 8'hec;
		memory[16'h1d94] <= 8'h14;
		memory[16'h1d95] <= 8'h3d;
		memory[16'h1d96] <= 8'hcf;
		memory[16'h1d97] <= 8'h75;
		memory[16'h1d98] <= 8'h9b;
		memory[16'h1d99] <= 8'h31;
		memory[16'h1d9a] <= 8'h0;
		memory[16'h1d9b] <= 8'h56;
		memory[16'h1d9c] <= 8'h81;
		memory[16'h1d9d] <= 8'h4f;
		memory[16'h1d9e] <= 8'h75;
		memory[16'h1d9f] <= 8'h57;
		memory[16'h1da0] <= 8'h13;
		memory[16'h1da1] <= 8'h38;
		memory[16'h1da2] <= 8'h7e;
		memory[16'h1da3] <= 8'h34;
		memory[16'h1da4] <= 8'h60;
		memory[16'h1da5] <= 8'h53;
		memory[16'h1da6] <= 8'h8c;
		memory[16'h1da7] <= 8'h30;
		memory[16'h1da8] <= 8'h12;
		memory[16'h1da9] <= 8'h34;
		memory[16'h1daa] <= 8'hbd;
		memory[16'h1dab] <= 8'he6;
		memory[16'h1dac] <= 8'h5f;
		memory[16'h1dad] <= 8'h24;
		memory[16'h1dae] <= 8'hbc;
		memory[16'h1daf] <= 8'h62;
		memory[16'h1db0] <= 8'hfd;
		memory[16'h1db1] <= 8'h62;
		memory[16'h1db2] <= 8'h4e;
		memory[16'h1db3] <= 8'h11;
		memory[16'h1db4] <= 8'h9f;
		memory[16'h1db5] <= 8'h1e;
		memory[16'h1db6] <= 8'h86;
		memory[16'h1db7] <= 8'h3b;
		memory[16'h1db8] <= 8'h4f;
		memory[16'h1db9] <= 8'h86;
		memory[16'h1dba] <= 8'h91;
		memory[16'h1dbb] <= 8'hd0;
		memory[16'h1dbc] <= 8'hd6;
		memory[16'h1dbd] <= 8'h6;
		memory[16'h1dbe] <= 8'h27;
		memory[16'h1dbf] <= 8'he9;
		memory[16'h1dc0] <= 8'h3e;
		memory[16'h1dc1] <= 8'ha5;
		memory[16'h1dc2] <= 8'h1e;
		memory[16'h1dc3] <= 8'h9f;
		memory[16'h1dc4] <= 8'hf8;
		memory[16'h1dc5] <= 8'haa;
		memory[16'h1dc6] <= 8'hcf;
		memory[16'h1dc7] <= 8'hb;
		memory[16'h1dc8] <= 8'hde;
		memory[16'h1dc9] <= 8'h8c;
		memory[16'h1dca] <= 8'hf1;
		memory[16'h1dcb] <= 8'h3e;
		memory[16'h1dcc] <= 8'hb0;
		memory[16'h1dcd] <= 8'hae;
		memory[16'h1dce] <= 8'ha0;
		memory[16'h1dcf] <= 8'had;
		memory[16'h1dd0] <= 8'h10;
		memory[16'h1dd1] <= 8'hee;
		memory[16'h1dd2] <= 8'hbf;
		memory[16'h1dd3] <= 8'haf;
		memory[16'h1dd4] <= 8'hc;
		memory[16'h1dd5] <= 8'h45;
		memory[16'h1dd6] <= 8'hea;
		memory[16'h1dd7] <= 8'h5b;
		memory[16'h1dd8] <= 8'hcc;
		memory[16'h1dd9] <= 8'h7b;
		memory[16'h1dda] <= 8'h2b;
		memory[16'h1ddb] <= 8'ha2;
		memory[16'h1ddc] <= 8'h81;
		memory[16'h1ddd] <= 8'h53;
		memory[16'h1dde] <= 8'h8b;
		memory[16'h1ddf] <= 8'hc0;
		memory[16'h1de0] <= 8'hf8;
		memory[16'h1de1] <= 8'ha9;
		memory[16'h1de2] <= 8'h5f;
		memory[16'h1de3] <= 8'hf1;
		memory[16'h1de4] <= 8'h54;
		memory[16'h1de5] <= 8'h2e;
		memory[16'h1de6] <= 8'hfc;
		memory[16'h1de7] <= 8'h32;
		memory[16'h1de8] <= 8'hbb;
		memory[16'h1de9] <= 8'hed;
		memory[16'h1dea] <= 8'h70;
		memory[16'h1deb] <= 8'h6b;
		memory[16'h1dec] <= 8'h9b;
		memory[16'h1ded] <= 8'h10;
		memory[16'h1dee] <= 8'h19;
		memory[16'h1def] <= 8'hab;
		memory[16'h1df0] <= 8'hff;
		memory[16'h1df1] <= 8'hd8;
		memory[16'h1df2] <= 8'h5b;
		memory[16'h1df3] <= 8'hb;
		memory[16'h1df4] <= 8'h1d;
		memory[16'h1df5] <= 8'h45;
		memory[16'h1df6] <= 8'h67;
		memory[16'h1df7] <= 8'he9;
		memory[16'h1df8] <= 8'hc1;
		memory[16'h1df9] <= 8'h92;
		memory[16'h1dfa] <= 8'h8b;
		memory[16'h1dfb] <= 8'h42;
		memory[16'h1dfc] <= 8'he5;
		memory[16'h1dfd] <= 8'h17;
		memory[16'h1dfe] <= 8'h2;
		memory[16'h1dff] <= 8'hde;
		memory[16'h1e00] <= 8'hc0;
		memory[16'h1e01] <= 8'h61;
		memory[16'h1e02] <= 8'hcf;
		memory[16'h1e03] <= 8'h14;
		memory[16'h1e04] <= 8'h90;
		memory[16'h1e05] <= 8'hcb;
		memory[16'h1e06] <= 8'h47;
		memory[16'h1e07] <= 8'h4b;
		memory[16'h1e08] <= 8'hb8;
		memory[16'h1e09] <= 8'hb7;
		memory[16'h1e0a] <= 8'hb6;
		memory[16'h1e0b] <= 8'h54;
		memory[16'h1e0c] <= 8'hc8;
		memory[16'h1e0d] <= 8'hcf;
		memory[16'h1e0e] <= 8'hff;
		memory[16'h1e0f] <= 8'hc7;
		memory[16'h1e10] <= 8'ha7;
		memory[16'h1e11] <= 8'h5a;
		memory[16'h1e12] <= 8'hd2;
		memory[16'h1e13] <= 8'hc5;
		memory[16'h1e14] <= 8'ha0;
		memory[16'h1e15] <= 8'h39;
		memory[16'h1e16] <= 8'hae;
		memory[16'h1e17] <= 8'h61;
		memory[16'h1e18] <= 8'hcc;
		memory[16'h1e19] <= 8'h3a;
		memory[16'h1e1a] <= 8'ha3;
		memory[16'h1e1b] <= 8'hb1;
		memory[16'h1e1c] <= 8'h51;
		memory[16'h1e1d] <= 8'ha6;
		memory[16'h1e1e] <= 8'h8f;
		memory[16'h1e1f] <= 8'h11;
		memory[16'h1e20] <= 8'h7;
		memory[16'h1e21] <= 8'h5e;
		memory[16'h1e22] <= 8'h26;
		memory[16'h1e23] <= 8'h97;
		memory[16'h1e24] <= 8'h29;
		memory[16'h1e25] <= 8'h6d;
		memory[16'h1e26] <= 8'he2;
		memory[16'h1e27] <= 8'he2;
		memory[16'h1e28] <= 8'h24;
		memory[16'h1e29] <= 8'h99;
		memory[16'h1e2a] <= 8'h36;
		memory[16'h1e2b] <= 8'hec;
		memory[16'h1e2c] <= 8'h68;
		memory[16'h1e2d] <= 8'h35;
		memory[16'h1e2e] <= 8'hb3;
		memory[16'h1e2f] <= 8'h10;
		memory[16'h1e30] <= 8'h90;
		memory[16'h1e31] <= 8'h86;
		memory[16'h1e32] <= 8'hd5;
		memory[16'h1e33] <= 8'h30;
		memory[16'h1e34] <= 8'hbf;
		memory[16'h1e35] <= 8'h83;
		memory[16'h1e36] <= 8'h91;
		memory[16'h1e37] <= 8'h8b;
		memory[16'h1e38] <= 8'hbd;
		memory[16'h1e39] <= 8'h34;
		memory[16'h1e3a] <= 8'h3d;
		memory[16'h1e3b] <= 8'he;
		memory[16'h1e3c] <= 8'hda;
		memory[16'h1e3d] <= 8'hcc;
		memory[16'h1e3e] <= 8'h20;
		memory[16'h1e3f] <= 8'he2;
		memory[16'h1e40] <= 8'h2b;
		memory[16'h1e41] <= 8'h46;
		memory[16'h1e42] <= 8'h79;
		memory[16'h1e43] <= 8'h54;
		memory[16'h1e44] <= 8'hb3;
		memory[16'h1e45] <= 8'h5c;
		memory[16'h1e46] <= 8'h36;
		memory[16'h1e47] <= 8'hd7;
		memory[16'h1e48] <= 8'hf5;
		memory[16'h1e49] <= 8'h6c;
		memory[16'h1e4a] <= 8'hc4;
		memory[16'h1e4b] <= 8'h5d;
		memory[16'h1e4c] <= 8'ha2;
		memory[16'h1e4d] <= 8'h77;
		memory[16'h1e4e] <= 8'h6d;
		memory[16'h1e4f] <= 8'h32;
		memory[16'h1e50] <= 8'hfd;
		memory[16'h1e51] <= 8'h42;
		memory[16'h1e52] <= 8'h62;
		memory[16'h1e53] <= 8'hbd;
		memory[16'h1e54] <= 8'hc6;
		memory[16'h1e55] <= 8'hf3;
		memory[16'h1e56] <= 8'h48;
		memory[16'h1e57] <= 8'h83;
		memory[16'h1e58] <= 8'h27;
		memory[16'h1e59] <= 8'h85;
		memory[16'h1e5a] <= 8'h92;
		memory[16'h1e5b] <= 8'h2;
		memory[16'h1e5c] <= 8'h52;
		memory[16'h1e5d] <= 8'hb2;
		memory[16'h1e5e] <= 8'he4;
		memory[16'h1e5f] <= 8'h7d;
		memory[16'h1e60] <= 8'hf8;
		memory[16'h1e61] <= 8'h5d;
		memory[16'h1e62] <= 8'hd1;
		memory[16'h1e63] <= 8'hab;
		memory[16'h1e64] <= 8'hb9;
		memory[16'h1e65] <= 8'h8;
		memory[16'h1e66] <= 8'h82;
		memory[16'h1e67] <= 8'hae;
		memory[16'h1e68] <= 8'h74;
		memory[16'h1e69] <= 8'h46;
		memory[16'h1e6a] <= 8'hc;
		memory[16'h1e6b] <= 8'h16;
		memory[16'h1e6c] <= 8'hbe;
		memory[16'h1e6d] <= 8'h79;
		memory[16'h1e6e] <= 8'h48;
		memory[16'h1e6f] <= 8'hbb;
		memory[16'h1e70] <= 8'hbc;
		memory[16'h1e71] <= 8'haa;
		memory[16'h1e72] <= 8'h78;
		memory[16'h1e73] <= 8'h82;
		memory[16'h1e74] <= 8'h9d;
		memory[16'h1e75] <= 8'hc1;
		memory[16'h1e76] <= 8'h5;
		memory[16'h1e77] <= 8'hc5;
		memory[16'h1e78] <= 8'h46;
		memory[16'h1e79] <= 8'h97;
		memory[16'h1e7a] <= 8'hc7;
		memory[16'h1e7b] <= 8'h98;
		memory[16'h1e7c] <= 8'h49;
		memory[16'h1e7d] <= 8'hab;
		memory[16'h1e7e] <= 8'h15;
		memory[16'h1e7f] <= 8'h41;
		memory[16'h1e80] <= 8'h8;
		memory[16'h1e81] <= 8'he7;
		memory[16'h1e82] <= 8'hec;
		memory[16'h1e83] <= 8'hc2;
		memory[16'h1e84] <= 8'hef;
		memory[16'h1e85] <= 8'h6f;
		memory[16'h1e86] <= 8'h70;
		memory[16'h1e87] <= 8'h63;
		memory[16'h1e88] <= 8'hb5;
		memory[16'h1e89] <= 8'h7c;
		memory[16'h1e8a] <= 8'h7a;
		memory[16'h1e8b] <= 8'h73;
		memory[16'h1e8c] <= 8'hf6;
		memory[16'h1e8d] <= 8'hc2;
		memory[16'h1e8e] <= 8'h2f;
		memory[16'h1e8f] <= 8'hb2;
		memory[16'h1e90] <= 8'h6d;
		memory[16'h1e91] <= 8'ha7;
		memory[16'h1e92] <= 8'h34;
		memory[16'h1e93] <= 8'ha;
		memory[16'h1e94] <= 8'h68;
		memory[16'h1e95] <= 8'h39;
		memory[16'h1e96] <= 8'hcf;
		memory[16'h1e97] <= 8'haf;
		memory[16'h1e98] <= 8'hd1;
		memory[16'h1e99] <= 8'h96;
		memory[16'h1e9a] <= 8'h47;
		memory[16'h1e9b] <= 8'h1a;
		memory[16'h1e9c] <= 8'h41;
		memory[16'h1e9d] <= 8'h5d;
		memory[16'h1e9e] <= 8'h5c;
		memory[16'h1e9f] <= 8'h4a;
		memory[16'h1ea0] <= 8'h44;
		memory[16'h1ea1] <= 8'h48;
		memory[16'h1ea2] <= 8'hc;
		memory[16'h1ea3] <= 8'h33;
		memory[16'h1ea4] <= 8'hb7;
		memory[16'h1ea5] <= 8'h7c;
		memory[16'h1ea6] <= 8'h96;
		memory[16'h1ea7] <= 8'h6d;
		memory[16'h1ea8] <= 8'hf9;
		memory[16'h1ea9] <= 8'h10;
		memory[16'h1eaa] <= 8'he0;
		memory[16'h1eab] <= 8'hef;
		memory[16'h1eac] <= 8'hd3;
		memory[16'h1ead] <= 8'hf;
		memory[16'h1eae] <= 8'ha1;
		memory[16'h1eaf] <= 8'h40;
		memory[16'h1eb0] <= 8'hb7;
		memory[16'h1eb1] <= 8'hd5;
		memory[16'h1eb2] <= 8'h4a;
		memory[16'h1eb3] <= 8'h1f;
		memory[16'h1eb4] <= 8'he;
		memory[16'h1eb5] <= 8'h1a;
		memory[16'h1eb6] <= 8'hce;
		memory[16'h1eb7] <= 8'hdf;
		memory[16'h1eb8] <= 8'hb0;
		memory[16'h1eb9] <= 8'h16;
		memory[16'h1eba] <= 8'hfa;
		memory[16'h1ebb] <= 8'hf2;
		memory[16'h1ebc] <= 8'h73;
		memory[16'h1ebd] <= 8'h56;
		memory[16'h1ebe] <= 8'h3c;
		memory[16'h1ebf] <= 8'hb7;
		memory[16'h1ec0] <= 8'h9e;
		memory[16'h1ec1] <= 8'h48;
		memory[16'h1ec2] <= 8'hea;
		memory[16'h1ec3] <= 8'h56;
		memory[16'h1ec4] <= 8'hc4;
		memory[16'h1ec5] <= 8'h80;
		memory[16'h1ec6] <= 8'hc3;
		memory[16'h1ec7] <= 8'hbd;
		memory[16'h1ec8] <= 8'h91;
		memory[16'h1ec9] <= 8'ha3;
		memory[16'h1eca] <= 8'hac;
		memory[16'h1ecb] <= 8'h64;
		memory[16'h1ecc] <= 8'hb3;
		memory[16'h1ecd] <= 8'h4d;
		memory[16'h1ece] <= 8'ha4;
		memory[16'h1ecf] <= 8'h6a;
		memory[16'h1ed0] <= 8'h22;
		memory[16'h1ed1] <= 8'hee;
		memory[16'h1ed2] <= 8'h89;
		memory[16'h1ed3] <= 8'h31;
		memory[16'h1ed4] <= 8'h8;
		memory[16'h1ed5] <= 8'h58;
		memory[16'h1ed6] <= 8'h10;
		memory[16'h1ed7] <= 8'hb9;
		memory[16'h1ed8] <= 8'h6e;
		memory[16'h1ed9] <= 8'ha;
		memory[16'h1eda] <= 8'hab;
		memory[16'h1edb] <= 8'he1;
		memory[16'h1edc] <= 8'h60;
		memory[16'h1edd] <= 8'he7;
		memory[16'h1ede] <= 8'h98;
		memory[16'h1edf] <= 8'hff;
		memory[16'h1ee0] <= 8'h2f;
		memory[16'h1ee1] <= 8'h82;
		memory[16'h1ee2] <= 8'h55;
		memory[16'h1ee3] <= 8'hf3;
		memory[16'h1ee4] <= 8'h2;
		memory[16'h1ee5] <= 8'h18;
		memory[16'h1ee6] <= 8'hb1;
		memory[16'h1ee7] <= 8'h93;
		memory[16'h1ee8] <= 8'hbb;
		memory[16'h1ee9] <= 8'h5d;
		memory[16'h1eea] <= 8'hf7;
		memory[16'h1eeb] <= 8'h6e;
		memory[16'h1eec] <= 8'hab;
		memory[16'h1eed] <= 8'h9b;
		memory[16'h1eee] <= 8'hd8;
		memory[16'h1eef] <= 8'hcd;
		memory[16'h1ef0] <= 8'h8a;
		memory[16'h1ef1] <= 8'h62;
		memory[16'h1ef2] <= 8'hfe;
		memory[16'h1ef3] <= 8'h92;
		memory[16'h1ef4] <= 8'hba;
		memory[16'h1ef5] <= 8'hf;
		memory[16'h1ef6] <= 8'h4b;
		memory[16'h1ef7] <= 8'h28;
		memory[16'h1ef8] <= 8'h19;
		memory[16'h1ef9] <= 8'hf6;
		memory[16'h1efa] <= 8'h9;
		memory[16'h1efb] <= 8'h7a;
		memory[16'h1efc] <= 8'hdd;
		memory[16'h1efd] <= 8'ha1;
		memory[16'h1efe] <= 8'h79;
		memory[16'h1eff] <= 8'hc;
		memory[16'h1f00] <= 8'h23;
		memory[16'h1f01] <= 8'hce;
		memory[16'h1f02] <= 8'h0;
		memory[16'h1f03] <= 8'h25;
		memory[16'h1f04] <= 8'he6;
		memory[16'h1f05] <= 8'hb1;
		memory[16'h1f06] <= 8'hb9;
		memory[16'h1f07] <= 8'ha1;
		memory[16'h1f08] <= 8'he;
		memory[16'h1f09] <= 8'hb0;
		memory[16'h1f0a] <= 8'h10;
		memory[16'h1f0b] <= 8'hb9;
		memory[16'h1f0c] <= 8'h4c;
		memory[16'h1f0d] <= 8'he8;
		memory[16'h1f0e] <= 8'h87;
		memory[16'h1f0f] <= 8'hd6;
		memory[16'h1f10] <= 8'h4a;
		memory[16'h1f11] <= 8'h85;
		memory[16'h1f12] <= 8'h68;
		memory[16'h1f13] <= 8'h4;
		memory[16'h1f14] <= 8'h94;
		memory[16'h1f15] <= 8'hb4;
		memory[16'h1f16] <= 8'h2c;
		memory[16'h1f17] <= 8'hae;
		memory[16'h1f18] <= 8'haa;
		memory[16'h1f19] <= 8'h35;
		memory[16'h1f1a] <= 8'h28;
		memory[16'h1f1b] <= 8'h88;
		memory[16'h1f1c] <= 8'hd6;
		memory[16'h1f1d] <= 8'ha1;
		memory[16'h1f1e] <= 8'h94;
		memory[16'h1f1f] <= 8'hf9;
		memory[16'h1f20] <= 8'h6f;
		memory[16'h1f21] <= 8'h94;
		memory[16'h1f22] <= 8'h1f;
		memory[16'h1f23] <= 8'h55;
		memory[16'h1f24] <= 8'h45;
		memory[16'h1f25] <= 8'hd8;
		memory[16'h1f26] <= 8'hf6;
		memory[16'h1f27] <= 8'h54;
		memory[16'h1f28] <= 8'h88;
		memory[16'h1f29] <= 8'h6;
		memory[16'h1f2a] <= 8'hd;
		memory[16'h1f2b] <= 8'hd4;
		memory[16'h1f2c] <= 8'hef;
		memory[16'h1f2d] <= 8'h94;
		memory[16'h1f2e] <= 8'haa;
		memory[16'h1f2f] <= 8'h39;
		memory[16'h1f30] <= 8'h1a;
		memory[16'h1f31] <= 8'h13;
		memory[16'h1f32] <= 8'h3e;
		memory[16'h1f33] <= 8'hae;
		memory[16'h1f34] <= 8'hc7;
		memory[16'h1f35] <= 8'h6a;
		memory[16'h1f36] <= 8'h5c;
		memory[16'h1f37] <= 8'h71;
		memory[16'h1f38] <= 8'ha0;
		memory[16'h1f39] <= 8'h84;
		memory[16'h1f3a] <= 8'hf9;
		memory[16'h1f3b] <= 8'h76;
		memory[16'h1f3c] <= 8'h25;
		memory[16'h1f3d] <= 8'h8e;
		memory[16'h1f3e] <= 8'h70;
		memory[16'h1f3f] <= 8'h94;
		memory[16'h1f40] <= 8'h22;
		memory[16'h1f41] <= 8'h8f;
		memory[16'h1f42] <= 8'he9;
		memory[16'h1f43] <= 8'h68;
		memory[16'h1f44] <= 8'h67;
		memory[16'h1f45] <= 8'he0;
		memory[16'h1f46] <= 8'hbc;
		memory[16'h1f47] <= 8'hef;
		memory[16'h1f48] <= 8'he6;
		memory[16'h1f49] <= 8'hc9;
		memory[16'h1f4a] <= 8'hc4;
		memory[16'h1f4b] <= 8'hd5;
		memory[16'h1f4c] <= 8'h5e;
		memory[16'h1f4d] <= 8'h6e;
		memory[16'h1f4e] <= 8'hf;
		memory[16'h1f4f] <= 8'h78;
		memory[16'h1f50] <= 8'h81;
		memory[16'h1f51] <= 8'h4d;
		memory[16'h1f52] <= 8'h26;
		memory[16'h1f53] <= 8'h48;
		memory[16'h1f54] <= 8'hb7;
		memory[16'h1f55] <= 8'h83;
		memory[16'h1f56] <= 8'hba;
		memory[16'h1f57] <= 8'h57;
		memory[16'h1f58] <= 8'h7;
		memory[16'h1f59] <= 8'hb3;
		memory[16'h1f5a] <= 8'hce;
		memory[16'h1f5b] <= 8'h2d;
		memory[16'h1f5c] <= 8'h41;
		memory[16'h1f5d] <= 8'h3e;
		memory[16'h1f5e] <= 8'hc1;
		memory[16'h1f5f] <= 8'h64;
		memory[16'h1f60] <= 8'hcd;
		memory[16'h1f61] <= 8'hab;
		memory[16'h1f62] <= 8'hcc;
		memory[16'h1f63] <= 8'h34;
		memory[16'h1f64] <= 8'h8b;
		memory[16'h1f65] <= 8'h88;
		memory[16'h1f66] <= 8'h23;
		memory[16'h1f67] <= 8'h71;
		memory[16'h1f68] <= 8'h51;
		memory[16'h1f69] <= 8'he7;
		memory[16'h1f6a] <= 8'h47;
		memory[16'h1f6b] <= 8'haf;
		memory[16'h1f6c] <= 8'h56;
		memory[16'h1f6d] <= 8'h56;
		memory[16'h1f6e] <= 8'h27;
		memory[16'h1f6f] <= 8'hd7;
		memory[16'h1f70] <= 8'ha3;
		memory[16'h1f71] <= 8'h4e;
		memory[16'h1f72] <= 8'h20;
		memory[16'h1f73] <= 8'h5a;
		memory[16'h1f74] <= 8'hd1;
		memory[16'h1f75] <= 8'hda;
		memory[16'h1f76] <= 8'hb2;
		memory[16'h1f77] <= 8'hd8;
		memory[16'h1f78] <= 8'h8d;
		memory[16'h1f79] <= 8'h80;
		memory[16'h1f7a] <= 8'h5;
		memory[16'h1f7b] <= 8'hcf;
		memory[16'h1f7c] <= 8'hbe;
		memory[16'h1f7d] <= 8'hc7;
		memory[16'h1f7e] <= 8'h33;
		memory[16'h1f7f] <= 8'h8b;
		memory[16'h1f80] <= 8'h72;
		memory[16'h1f81] <= 8'hff;
		memory[16'h1f82] <= 8'hbf;
		memory[16'h1f83] <= 8'hfd;
		memory[16'h1f84] <= 8'h87;
		memory[16'h1f85] <= 8'he2;
		memory[16'h1f86] <= 8'h6e;
		memory[16'h1f87] <= 8'hd8;
		memory[16'h1f88] <= 8'hca;
		memory[16'h1f89] <= 8'hb5;
		memory[16'h1f8a] <= 8'h88;
		memory[16'h1f8b] <= 8'h20;
		memory[16'h1f8c] <= 8'hb;
		memory[16'h1f8d] <= 8'haf;
		memory[16'h1f8e] <= 8'hf7;
		memory[16'h1f8f] <= 8'hae;
		memory[16'h1f90] <= 8'hfd;
		memory[16'h1f91] <= 8'h17;
		memory[16'h1f92] <= 8'h9;
		memory[16'h1f93] <= 8'hce;
		memory[16'h1f94] <= 8'hf1;
		memory[16'h1f95] <= 8'hbb;
		memory[16'h1f96] <= 8'ha7;
		memory[16'h1f97] <= 8'h7f;
		memory[16'h1f98] <= 8'h3b;
		memory[16'h1f99] <= 8'hac;
		memory[16'h1f9a] <= 8'h4e;
		memory[16'h1f9b] <= 8'hf9;
		memory[16'h1f9c] <= 8'h73;
		memory[16'h1f9d] <= 8'h81;
		memory[16'h1f9e] <= 8'h84;
		memory[16'h1f9f] <= 8'he5;
		memory[16'h1fa0] <= 8'h80;
		memory[16'h1fa1] <= 8'h43;
		memory[16'h1fa2] <= 8'he2;
		memory[16'h1fa3] <= 8'h7;
		memory[16'h1fa4] <= 8'h25;
		memory[16'h1fa5] <= 8'h51;
		memory[16'h1fa6] <= 8'hdf;
		memory[16'h1fa7] <= 8'hef;
		memory[16'h1fa8] <= 8'h6;
		memory[16'h1fa9] <= 8'h67;
		memory[16'h1faa] <= 8'hf;
		memory[16'h1fab] <= 8'h12;
		memory[16'h1fac] <= 8'h17;
		memory[16'h1fad] <= 8'h7;
		memory[16'h1fae] <= 8'hc0;
		memory[16'h1faf] <= 8'h14;
		memory[16'h1fb0] <= 8'h1e;
		memory[16'h1fb1] <= 8'hc9;
		memory[16'h1fb2] <= 8'he3;
		memory[16'h1fb3] <= 8'h10;
		memory[16'h1fb4] <= 8'h84;
		memory[16'h1fb5] <= 8'h8a;
		memory[16'h1fb6] <= 8'h8f;
		memory[16'h1fb7] <= 8'hbf;
		memory[16'h1fb8] <= 8'h36;
		memory[16'h1fb9] <= 8'hdd;
		memory[16'h1fba] <= 8'hb8;
		memory[16'h1fbb] <= 8'haa;
		memory[16'h1fbc] <= 8'h5e;
		memory[16'h1fbd] <= 8'h3c;
		memory[16'h1fbe] <= 8'h8f;
		memory[16'h1fbf] <= 8'hde;
		memory[16'h1fc0] <= 8'h7f;
		memory[16'h1fc1] <= 8'h72;
		memory[16'h1fc2] <= 8'he5;
		memory[16'h1fc3] <= 8'ha5;
		memory[16'h1fc4] <= 8'hc3;
		memory[16'h1fc5] <= 8'hc4;
		memory[16'h1fc6] <= 8'h94;
		memory[16'h1fc7] <= 8'hc9;
		memory[16'h1fc8] <= 8'h2c;
		memory[16'h1fc9] <= 8'ha4;
		memory[16'h1fca] <= 8'hdb;
		memory[16'h1fcb] <= 8'h43;
		memory[16'h1fcc] <= 8'hab;
		memory[16'h1fcd] <= 8'h9c;
		memory[16'h1fce] <= 8'h57;
		memory[16'h1fcf] <= 8'hc9;
		memory[16'h1fd0] <= 8'h65;
		memory[16'h1fd1] <= 8'h3a;
		memory[16'h1fd2] <= 8'hd9;
		memory[16'h1fd3] <= 8'hea;
		memory[16'h1fd4] <= 8'hc4;
		memory[16'h1fd5] <= 8'h68;
		memory[16'h1fd6] <= 8'ha9;
		memory[16'h1fd7] <= 8'hfb;
		memory[16'h1fd8] <= 8'h45;
		memory[16'h1fd9] <= 8'h62;
		memory[16'h1fda] <= 8'ha5;
		memory[16'h1fdb] <= 8'ha3;
		memory[16'h1fdc] <= 8'h9e;
		memory[16'h1fdd] <= 8'h34;
		memory[16'h1fde] <= 8'h81;
		memory[16'h1fdf] <= 8'h1e;
		memory[16'h1fe0] <= 8'ha6;
		memory[16'h1fe1] <= 8'h66;
		memory[16'h1fe2] <= 8'hc3;
		memory[16'h1fe3] <= 8'h69;
		memory[16'h1fe4] <= 8'h2b;
		memory[16'h1fe5] <= 8'h57;
		memory[16'h1fe6] <= 8'h33;
		memory[16'h1fe7] <= 8'h57;
		memory[16'h1fe8] <= 8'hfb;
		memory[16'h1fe9] <= 8'he;
		memory[16'h1fea] <= 8'h9a;
		memory[16'h1feb] <= 8'ha6;
		memory[16'h1fec] <= 8'haa;
		memory[16'h1fed] <= 8'hf1;
		memory[16'h1fee] <= 8'h70;
		memory[16'h1fef] <= 8'h10;
		memory[16'h1ff0] <= 8'h2c;
		memory[16'h1ff1] <= 8'h49;
		memory[16'h1ff2] <= 8'hfa;
		memory[16'h1ff3] <= 8'hf0;
		memory[16'h1ff4] <= 8'hb2;
		memory[16'h1ff5] <= 8'ha3;
		memory[16'h1ff6] <= 8'heb;
		memory[16'h1ff7] <= 8'hf7;
		memory[16'h1ff8] <= 8'h5;
		memory[16'h1ff9] <= 8'h90;
		memory[16'h1ffa] <= 8'h9b;
		memory[16'h1ffb] <= 8'ha4;
		memory[16'h1ffc] <= 8'hc5;
		memory[16'h1ffd] <= 8'h1c;
		memory[16'h1ffe] <= 8'hc2;
		memory[16'h1fff] <= 8'h6b;
		memory[16'h2000] <= 8'h83;
		memory[16'h2001] <= 8'h85;
		memory[16'h2002] <= 8'hd5;
		memory[16'h2003] <= 8'hae;
		memory[16'h2004] <= 8'hdc;
		memory[16'h2005] <= 8'h8;
		memory[16'h2006] <= 8'h5;
		memory[16'h2007] <= 8'hd8;
		memory[16'h2008] <= 8'h16;
		memory[16'h2009] <= 8'h9f;
		memory[16'h200a] <= 8'h7e;
		memory[16'h200b] <= 8'hc1;
		memory[16'h200c] <= 8'h90;
		memory[16'h200d] <= 8'hee;
		memory[16'h200e] <= 8'hd1;
		memory[16'h200f] <= 8'hbc;
		memory[16'h2010] <= 8'h38;
		memory[16'h2011] <= 8'hcb;
		memory[16'h2012] <= 8'had;
		memory[16'h2013] <= 8'hea;
		memory[16'h2014] <= 8'h6e;
		memory[16'h2015] <= 8'h98;
		memory[16'h2016] <= 8'he1;
		memory[16'h2017] <= 8'h74;
		memory[16'h2018] <= 8'h29;
		memory[16'h2019] <= 8'h7c;
		memory[16'h201a] <= 8'h18;
		memory[16'h201b] <= 8'hee;
		memory[16'h201c] <= 8'h99;
		memory[16'h201d] <= 8'hda;
		memory[16'h201e] <= 8'h59;
		memory[16'h201f] <= 8'h1c;
		memory[16'h2020] <= 8'h5f;
		memory[16'h2021] <= 8'h2e;
		memory[16'h2022] <= 8'hca;
		memory[16'h2023] <= 8'h3b;
		memory[16'h2024] <= 8'h36;
		memory[16'h2025] <= 8'hcf;
		memory[16'h2026] <= 8'h13;
		memory[16'h2027] <= 8'h4d;
		memory[16'h2028] <= 8'h6e;
		memory[16'h2029] <= 8'h92;
		memory[16'h202a] <= 8'he;
		memory[16'h202b] <= 8'hfe;
		memory[16'h202c] <= 8'h80;
		memory[16'h202d] <= 8'hdf;
		memory[16'h202e] <= 8'hbb;
		memory[16'h202f] <= 8'hb8;
		memory[16'h2030] <= 8'haa;
		memory[16'h2031] <= 8'h68;
		memory[16'h2032] <= 8'ha2;
		memory[16'h2033] <= 8'h18;
		memory[16'h2034] <= 8'h0;
		memory[16'h2035] <= 8'h84;
		memory[16'h2036] <= 8'h8c;
		memory[16'h2037] <= 8'h29;
		memory[16'h2038] <= 8'h0;
		memory[16'h2039] <= 8'ha4;
		memory[16'h203a] <= 8'h17;
		memory[16'h203b] <= 8'h99;
		memory[16'h203c] <= 8'h7e;
		memory[16'h203d] <= 8'h71;
		memory[16'h203e] <= 8'hb5;
		memory[16'h203f] <= 8'hdd;
		memory[16'h2040] <= 8'h9f;
		memory[16'h2041] <= 8'h7f;
		memory[16'h2042] <= 8'h19;
		memory[16'h2043] <= 8'hd6;
		memory[16'h2044] <= 8'h4e;
		memory[16'h2045] <= 8'h2c;
		memory[16'h2046] <= 8'h23;
		memory[16'h2047] <= 8'hbc;
		memory[16'h2048] <= 8'hbe;
		memory[16'h2049] <= 8'h31;
		memory[16'h204a] <= 8'hbb;
		memory[16'h204b] <= 8'h3f;
		memory[16'h204c] <= 8'h10;
		memory[16'h204d] <= 8'h76;
		memory[16'h204e] <= 8'hf7;
		memory[16'h204f] <= 8'hba;
		memory[16'h2050] <= 8'hde;
		memory[16'h2051] <= 8'h9a;
		memory[16'h2052] <= 8'hd2;
		memory[16'h2053] <= 8'hde;
		memory[16'h2054] <= 8'h1e;
		memory[16'h2055] <= 8'h5f;
		memory[16'h2056] <= 8'h8;
		memory[16'h2057] <= 8'h1e;
		memory[16'h2058] <= 8'h3;
		memory[16'h2059] <= 8'h1f;
		memory[16'h205a] <= 8'hb8;
		memory[16'h205b] <= 8'h82;
		memory[16'h205c] <= 8'h90;
		memory[16'h205d] <= 8'h6d;
		memory[16'h205e] <= 8'h5f;
		memory[16'h205f] <= 8'h30;
		memory[16'h2060] <= 8'hed;
		memory[16'h2061] <= 8'h78;
		memory[16'h2062] <= 8'h6;
		memory[16'h2063] <= 8'h3b;
		memory[16'h2064] <= 8'ha5;
		memory[16'h2065] <= 8'h29;
		memory[16'h2066] <= 8'hf8;
		memory[16'h2067] <= 8'h63;
		memory[16'h2068] <= 8'h5a;
		memory[16'h2069] <= 8'hb3;
		memory[16'h206a] <= 8'ha2;
		memory[16'h206b] <= 8'h6a;
		memory[16'h206c] <= 8'h29;
		memory[16'h206d] <= 8'h9a;
		memory[16'h206e] <= 8'h24;
		memory[16'h206f] <= 8'h7;
		memory[16'h2070] <= 8'h34;
		memory[16'h2071] <= 8'hf6;
		memory[16'h2072] <= 8'he5;
		memory[16'h2073] <= 8'h52;
		memory[16'h2074] <= 8'h55;
		memory[16'h2075] <= 8'hed;
		memory[16'h2076] <= 8'h70;
		memory[16'h2077] <= 8'h59;
		memory[16'h2078] <= 8'hd;
		memory[16'h2079] <= 8'h28;
		memory[16'h207a] <= 8'hdb;
		memory[16'h207b] <= 8'h9d;
		memory[16'h207c] <= 8'h96;
		memory[16'h207d] <= 8'h3a;
		memory[16'h207e] <= 8'hcd;
		memory[16'h207f] <= 8'h83;
		memory[16'h2080] <= 8'hb3;
		memory[16'h2081] <= 8'hd3;
		memory[16'h2082] <= 8'hbe;
		memory[16'h2083] <= 8'h58;
		memory[16'h2084] <= 8'hfc;
		memory[16'h2085] <= 8'hb6;
		memory[16'h2086] <= 8'hbb;
		memory[16'h2087] <= 8'h56;
		memory[16'h2088] <= 8'h69;
		memory[16'h2089] <= 8'h5e;
		memory[16'h208a] <= 8'hc0;
		memory[16'h208b] <= 8'h92;
		memory[16'h208c] <= 8'hf8;
		memory[16'h208d] <= 8'he4;
		memory[16'h208e] <= 8'h99;
		memory[16'h208f] <= 8'h2c;
		memory[16'h2090] <= 8'hdb;
		memory[16'h2091] <= 8'h7f;
		memory[16'h2092] <= 8'h7e;
		memory[16'h2093] <= 8'h30;
		memory[16'h2094] <= 8'h6c;
		memory[16'h2095] <= 8'hee;
		memory[16'h2096] <= 8'h89;
		memory[16'h2097] <= 8'h79;
		memory[16'h2098] <= 8'h17;
		memory[16'h2099] <= 8'h64;
		memory[16'h209a] <= 8'h17;
		memory[16'h209b] <= 8'had;
		memory[16'h209c] <= 8'h9f;
		memory[16'h209d] <= 8'he4;
		memory[16'h209e] <= 8'h30;
		memory[16'h209f] <= 8'h52;
		memory[16'h20a0] <= 8'hb8;
		memory[16'h20a1] <= 8'hee;
		memory[16'h20a2] <= 8'haa;
		memory[16'h20a3] <= 8'hb4;
		memory[16'h20a4] <= 8'ha5;
		memory[16'h20a5] <= 8'h65;
		memory[16'h20a6] <= 8'hb;
		memory[16'h20a7] <= 8'he;
		memory[16'h20a8] <= 8'hc3;
		memory[16'h20a9] <= 8'hcb;
		memory[16'h20aa] <= 8'ha1;
		memory[16'h20ab] <= 8'hbb;
		memory[16'h20ac] <= 8'hb0;
		memory[16'h20ad] <= 8'h3a;
		memory[16'h20ae] <= 8'he7;
		memory[16'h20af] <= 8'h8b;
		memory[16'h20b0] <= 8'hb9;
		memory[16'h20b1] <= 8'h65;
		memory[16'h20b2] <= 8'hbb;
		memory[16'h20b3] <= 8'h26;
		memory[16'h20b4] <= 8'h54;
		memory[16'h20b5] <= 8'h45;
		memory[16'h20b6] <= 8'h9f;
		memory[16'h20b7] <= 8'h6b;
		memory[16'h20b8] <= 8'ha9;
		memory[16'h20b9] <= 8'hb6;
		memory[16'h20ba] <= 8'h18;
		memory[16'h20bb] <= 8'h48;
		memory[16'h20bc] <= 8'h9b;
		memory[16'h20bd] <= 8'h48;
		memory[16'h20be] <= 8'h9a;
		memory[16'h20bf] <= 8'h53;
		memory[16'h20c0] <= 8'h36;
		memory[16'h20c1] <= 8'h44;
		memory[16'h20c2] <= 8'h7;
		memory[16'h20c3] <= 8'hdb;
		memory[16'h20c4] <= 8'haa;
		memory[16'h20c5] <= 8'h12;
		memory[16'h20c6] <= 8'hea;
		memory[16'h20c7] <= 8'h6d;
		memory[16'h20c8] <= 8'hde;
		memory[16'h20c9] <= 8'h8b;
		memory[16'h20ca] <= 8'h29;
		memory[16'h20cb] <= 8'h8e;
		memory[16'h20cc] <= 8'hc5;
		memory[16'h20cd] <= 8'h10;
		memory[16'h20ce] <= 8'h19;
		memory[16'h20cf] <= 8'h7f;
		memory[16'h20d0] <= 8'h76;
		memory[16'h20d1] <= 8'hd4;
		memory[16'h20d2] <= 8'ha5;
		memory[16'h20d3] <= 8'hca;
		memory[16'h20d4] <= 8'h19;
		memory[16'h20d5] <= 8'h44;
		memory[16'h20d6] <= 8'h35;
		memory[16'h20d7] <= 8'hc3;
		memory[16'h20d8] <= 8'hfb;
		memory[16'h20d9] <= 8'h4d;
		memory[16'h20da] <= 8'hb;
		memory[16'h20db] <= 8'h96;
		memory[16'h20dc] <= 8'h95;
		memory[16'h20dd] <= 8'ha6;
		memory[16'h20de] <= 8'he9;
		memory[16'h20df] <= 8'hcb;
		memory[16'h20e0] <= 8'hea;
		memory[16'h20e1] <= 8'hf0;
		memory[16'h20e2] <= 8'ha7;
		memory[16'h20e3] <= 8'h94;
		memory[16'h20e4] <= 8'h3;
		memory[16'h20e5] <= 8'h91;
		memory[16'h20e6] <= 8'h2;
		memory[16'h20e7] <= 8'he1;
		memory[16'h20e8] <= 8'h1c;
		memory[16'h20e9] <= 8'h2b;
		memory[16'h20ea] <= 8'h6f;
		memory[16'h20eb] <= 8'he1;
		memory[16'h20ec] <= 8'h3b;
		memory[16'h20ed] <= 8'h88;
		memory[16'h20ee] <= 8'h60;
		memory[16'h20ef] <= 8'hb1;
		memory[16'h20f0] <= 8'h5c;
		memory[16'h20f1] <= 8'h5;
		memory[16'h20f2] <= 8'h7b;
		memory[16'h20f3] <= 8'h76;
		memory[16'h20f4] <= 8'h4a;
		memory[16'h20f5] <= 8'hb0;
		memory[16'h20f6] <= 8'h39;
		memory[16'h20f7] <= 8'h45;
		memory[16'h20f8] <= 8'hfd;
		memory[16'h20f9] <= 8'h44;
		memory[16'h20fa] <= 8'hdb;
		memory[16'h20fb] <= 8'h92;
		memory[16'h20fc] <= 8'hea;
		memory[16'h20fd] <= 8'hc4;
		memory[16'h20fe] <= 8'h5e;
		memory[16'h20ff] <= 8'hd5;
		memory[16'h2100] <= 8'hb4;
		memory[16'h2101] <= 8'h5;
		memory[16'h2102] <= 8'h69;
		memory[16'h2103] <= 8'hb7;
		memory[16'h2104] <= 8'h96;
		memory[16'h2105] <= 8'h6b;
		memory[16'h2106] <= 8'h98;
		memory[16'h2107] <= 8'hb2;
		memory[16'h2108] <= 8'h96;
		memory[16'h2109] <= 8'h7;
		memory[16'h210a] <= 8'h93;
		memory[16'h210b] <= 8'hd2;
		memory[16'h210c] <= 8'h8f;
		memory[16'h210d] <= 8'hf4;
		memory[16'h210e] <= 8'h83;
		memory[16'h210f] <= 8'hec;
		memory[16'h2110] <= 8'hf9;
		memory[16'h2111] <= 8'hff;
		memory[16'h2112] <= 8'h62;
		memory[16'h2113] <= 8'h43;
		memory[16'h2114] <= 8'haf;
		memory[16'h2115] <= 8'h9b;
		memory[16'h2116] <= 8'h88;
		memory[16'h2117] <= 8'had;
		memory[16'h2118] <= 8'hdf;
		memory[16'h2119] <= 8'h63;
		memory[16'h211a] <= 8'h3f;
		memory[16'h211b] <= 8'hca;
		memory[16'h211c] <= 8'h27;
		memory[16'h211d] <= 8'h9d;
		memory[16'h211e] <= 8'h9f;
		memory[16'h211f] <= 8'hdc;
		memory[16'h2120] <= 8'ha2;
		memory[16'h2121] <= 8'h8;
		memory[16'h2122] <= 8'h93;
		memory[16'h2123] <= 8'h38;
		memory[16'h2124] <= 8'h74;
		memory[16'h2125] <= 8'h2c;
		memory[16'h2126] <= 8'hea;
		memory[16'h2127] <= 8'ha;
		memory[16'h2128] <= 8'h33;
		memory[16'h2129] <= 8'h7e;
		memory[16'h212a] <= 8'hdc;
		memory[16'h212b] <= 8'hc3;
		memory[16'h212c] <= 8'h72;
		memory[16'h212d] <= 8'h60;
		memory[16'h212e] <= 8'haf;
		memory[16'h212f] <= 8'h6b;
		memory[16'h2130] <= 8'h5f;
		memory[16'h2131] <= 8'h11;
		memory[16'h2132] <= 8'haf;
		memory[16'h2133] <= 8'he;
		memory[16'h2134] <= 8'hac;
		memory[16'h2135] <= 8'h37;
		memory[16'h2136] <= 8'hbb;
		memory[16'h2137] <= 8'h8b;
		memory[16'h2138] <= 8'h9b;
		memory[16'h2139] <= 8'hfb;
		memory[16'h213a] <= 8'h55;
		memory[16'h213b] <= 8'hc2;
		memory[16'h213c] <= 8'h98;
		memory[16'h213d] <= 8'hf4;
		memory[16'h213e] <= 8'h9e;
		memory[16'h213f] <= 8'h3b;
		memory[16'h2140] <= 8'hfd;
		memory[16'h2141] <= 8'h32;
		memory[16'h2142] <= 8'h73;
		memory[16'h2143] <= 8'h71;
		memory[16'h2144] <= 8'h5e;
		memory[16'h2145] <= 8'h5e;
		memory[16'h2146] <= 8'h7b;
		memory[16'h2147] <= 8'h91;
		memory[16'h2148] <= 8'hdc;
		memory[16'h2149] <= 8'h58;
		memory[16'h214a] <= 8'h54;
		memory[16'h214b] <= 8'h4e;
		memory[16'h214c] <= 8'hb8;
		memory[16'h214d] <= 8'h3;
		memory[16'h214e] <= 8'hb9;
		memory[16'h214f] <= 8'h17;
		memory[16'h2150] <= 8'h14;
		memory[16'h2151] <= 8'h68;
		memory[16'h2152] <= 8'h25;
		memory[16'h2153] <= 8'hc0;
		memory[16'h2154] <= 8'ha0;
		memory[16'h2155] <= 8'he1;
		memory[16'h2156] <= 8'h4c;
		memory[16'h2157] <= 8'h3b;
		memory[16'h2158] <= 8'hdc;
		memory[16'h2159] <= 8'ha1;
		memory[16'h215a] <= 8'hfd;
		memory[16'h215b] <= 8'h74;
		memory[16'h215c] <= 8'h96;
		memory[16'h215d] <= 8'h9c;
		memory[16'h215e] <= 8'haf;
		memory[16'h215f] <= 8'h93;
		memory[16'h2160] <= 8'hce;
		memory[16'h2161] <= 8'h23;
		memory[16'h2162] <= 8'h4;
		memory[16'h2163] <= 8'h2c;
		memory[16'h2164] <= 8'h81;
		memory[16'h2165] <= 8'h7f;
		memory[16'h2166] <= 8'hbd;
		memory[16'h2167] <= 8'h5d;
		memory[16'h2168] <= 8'hd7;
		memory[16'h2169] <= 8'h12;
		memory[16'h216a] <= 8'hab;
		memory[16'h216b] <= 8'h8f;
		memory[16'h216c] <= 8'h15;
		memory[16'h216d] <= 8'h64;
		memory[16'h216e] <= 8'ha6;
		memory[16'h216f] <= 8'h2a;
		memory[16'h2170] <= 8'hcd;
		memory[16'h2171] <= 8'hcc;
		memory[16'h2172] <= 8'hea;
		memory[16'h2173] <= 8'h6d;
		memory[16'h2174] <= 8'had;
		memory[16'h2175] <= 8'h36;
		memory[16'h2176] <= 8'ha8;
		memory[16'h2177] <= 8'h89;
		memory[16'h2178] <= 8'hd8;
		memory[16'h2179] <= 8'ha5;
		memory[16'h217a] <= 8'hfd;
		memory[16'h217b] <= 8'h6e;
		memory[16'h217c] <= 8'h41;
		memory[16'h217d] <= 8'had;
		memory[16'h217e] <= 8'h1;
		memory[16'h217f] <= 8'hf;
		memory[16'h2180] <= 8'hd0;
		memory[16'h2181] <= 8'h5;
		memory[16'h2182] <= 8'h3b;
		memory[16'h2183] <= 8'h51;
		memory[16'h2184] <= 8'h84;
		memory[16'h2185] <= 8'hf9;
		memory[16'h2186] <= 8'hae;
		memory[16'h2187] <= 8'h5c;
		memory[16'h2188] <= 8'hb;
		memory[16'h2189] <= 8'h59;
		memory[16'h218a] <= 8'heb;
		memory[16'h218b] <= 8'h20;
		memory[16'h218c] <= 8'hbd;
		memory[16'h218d] <= 8'h92;
		memory[16'h218e] <= 8'h4a;
		memory[16'h218f] <= 8'h8a;
		memory[16'h2190] <= 8'h5e;
		memory[16'h2191] <= 8'h35;
		memory[16'h2192] <= 8'hf7;
		memory[16'h2193] <= 8'hb;
		memory[16'h2194] <= 8'h6b;
		memory[16'h2195] <= 8'h9f;
		memory[16'h2196] <= 8'h94;
		memory[16'h2197] <= 8'h43;
		memory[16'h2198] <= 8'h45;
		memory[16'h2199] <= 8'h91;
		memory[16'h219a] <= 8'hb1;
		memory[16'h219b] <= 8'h86;
		memory[16'h219c] <= 8'h3e;
		memory[16'h219d] <= 8'hb2;
		memory[16'h219e] <= 8'h96;
		memory[16'h219f] <= 8'he;
		memory[16'h21a0] <= 8'hb7;
		memory[16'h21a1] <= 8'hd1;
		memory[16'h21a2] <= 8'h5f;
		memory[16'h21a3] <= 8'h3c;
		memory[16'h21a4] <= 8'hca;
		memory[16'h21a5] <= 8'hd;
		memory[16'h21a6] <= 8'h98;
		memory[16'h21a7] <= 8'hd5;
		memory[16'h21a8] <= 8'h66;
		memory[16'h21a9] <= 8'h83;
		memory[16'h21aa] <= 8'hf6;
		memory[16'h21ab] <= 8'h24;
		memory[16'h21ac] <= 8'h15;
		memory[16'h21ad] <= 8'h40;
		memory[16'h21ae] <= 8'hae;
		memory[16'h21af] <= 8'h73;
		memory[16'h21b0] <= 8'h75;
		memory[16'h21b1] <= 8'ha6;
		memory[16'h21b2] <= 8'h7e;
		memory[16'h21b3] <= 8'he1;
		memory[16'h21b4] <= 8'h45;
		memory[16'h21b5] <= 8'h12;
		memory[16'h21b6] <= 8'h24;
		memory[16'h21b7] <= 8'h8a;
		memory[16'h21b8] <= 8'ha4;
		memory[16'h21b9] <= 8'hd6;
		memory[16'h21ba] <= 8'h11;
		memory[16'h21bb] <= 8'he2;
		memory[16'h21bc] <= 8'h88;
		memory[16'h21bd] <= 8'ha7;
		memory[16'h21be] <= 8'hf1;
		memory[16'h21bf] <= 8'h40;
		memory[16'h21c0] <= 8'h78;
		memory[16'h21c1] <= 8'h50;
		memory[16'h21c2] <= 8'h7c;
		memory[16'h21c3] <= 8'h43;
		memory[16'h21c4] <= 8'h5e;
		memory[16'h21c5] <= 8'h14;
		memory[16'h21c6] <= 8'h18;
		memory[16'h21c7] <= 8'hc4;
		memory[16'h21c8] <= 8'h97;
		memory[16'h21c9] <= 8'he;
		memory[16'h21ca] <= 8'he8;
		memory[16'h21cb] <= 8'had;
		memory[16'h21cc] <= 8'h4f;
		memory[16'h21cd] <= 8'h97;
		memory[16'h21ce] <= 8'h20;
		memory[16'h21cf] <= 8'hc4;
		memory[16'h21d0] <= 8'h3d;
		memory[16'h21d1] <= 8'h9f;
		memory[16'h21d2] <= 8'ha5;
		memory[16'h21d3] <= 8'h82;
		memory[16'h21d4] <= 8'hb1;
		memory[16'h21d5] <= 8'hca;
		memory[16'h21d6] <= 8'hd;
		memory[16'h21d7] <= 8'h55;
		memory[16'h21d8] <= 8'ha0;
		memory[16'h21d9] <= 8'h1e;
		memory[16'h21da] <= 8'h38;
		memory[16'h21db] <= 8'h28;
		memory[16'h21dc] <= 8'hc5;
		memory[16'h21dd] <= 8'h29;
		memory[16'h21de] <= 8'h68;
		memory[16'h21df] <= 8'h3d;
		memory[16'h21e0] <= 8'h79;
		memory[16'h21e1] <= 8'he4;
		memory[16'h21e2] <= 8'h80;
		memory[16'h21e3] <= 8'hd7;
		memory[16'h21e4] <= 8'hf8;
		memory[16'h21e5] <= 8'h99;
		memory[16'h21e6] <= 8'h9c;
		memory[16'h21e7] <= 8'h90;
		memory[16'h21e8] <= 8'ha7;
		memory[16'h21e9] <= 8'h84;
		memory[16'h21ea] <= 8'h3d;
		memory[16'h21eb] <= 8'hf6;
		memory[16'h21ec] <= 8'h1b;
		memory[16'h21ed] <= 8'h5d;
		memory[16'h21ee] <= 8'hbb;
		memory[16'h21ef] <= 8'h58;
		memory[16'h21f0] <= 8'hfc;
		memory[16'h21f1] <= 8'h60;
		memory[16'h21f2] <= 8'hdb;
		memory[16'h21f3] <= 8'hae;
		memory[16'h21f4] <= 8'h2a;
		memory[16'h21f5] <= 8'he8;
		memory[16'h21f6] <= 8'h3;
		memory[16'h21f7] <= 8'hca;
		memory[16'h21f8] <= 8'h6;
		memory[16'h21f9] <= 8'h3b;
		memory[16'h21fa] <= 8'hf3;
		memory[16'h21fb] <= 8'hcb;
		memory[16'h21fc] <= 8'h64;
		memory[16'h21fd] <= 8'h5b;
		memory[16'h21fe] <= 8'h8;
		memory[16'h21ff] <= 8'hde;
		memory[16'h2200] <= 8'h40;
		memory[16'h2201] <= 8'h89;
		memory[16'h2202] <= 8'hb5;
		memory[16'h2203] <= 8'h38;
		memory[16'h2204] <= 8'h22;
		memory[16'h2205] <= 8'h51;
		memory[16'h2206] <= 8'hc8;
		memory[16'h2207] <= 8'hc9;
		memory[16'h2208] <= 8'hd6;
		memory[16'h2209] <= 8'h5;
		memory[16'h220a] <= 8'hc0;
		memory[16'h220b] <= 8'hf1;
		memory[16'h220c] <= 8'h63;
		memory[16'h220d] <= 8'h7b;
		memory[16'h220e] <= 8'h4a;
		memory[16'h220f] <= 8'h5f;
		memory[16'h2210] <= 8'hdb;
		memory[16'h2211] <= 8'h25;
		memory[16'h2212] <= 8'hd;
		memory[16'h2213] <= 8'h6;
		memory[16'h2214] <= 8'hd;
		memory[16'h2215] <= 8'h11;
		memory[16'h2216] <= 8'hd0;
		memory[16'h2217] <= 8'h13;
		memory[16'h2218] <= 8'h4c;
		memory[16'h2219] <= 8'hc3;
		memory[16'h221a] <= 8'hde;
		memory[16'h221b] <= 8'hb1;
		memory[16'h221c] <= 8'h1f;
		memory[16'h221d] <= 8'he6;
		memory[16'h221e] <= 8'h8f;
		memory[16'h221f] <= 8'h5f;
		memory[16'h2220] <= 8'h6f;
		memory[16'h2221] <= 8'h44;
		memory[16'h2222] <= 8'h97;
		memory[16'h2223] <= 8'h91;
		memory[16'h2224] <= 8'h96;
		memory[16'h2225] <= 8'h60;
		memory[16'h2226] <= 8'h5b;
		memory[16'h2227] <= 8'h6c;
		memory[16'h2228] <= 8'h65;
		memory[16'h2229] <= 8'h1b;
		memory[16'h222a] <= 8'h5d;
		memory[16'h222b] <= 8'hc8;
		memory[16'h222c] <= 8'h96;
		memory[16'h222d] <= 8'ha7;
		memory[16'h222e] <= 8'h28;
		memory[16'h222f] <= 8'h71;
		memory[16'h2230] <= 8'hcc;
		memory[16'h2231] <= 8'h35;
		memory[16'h2232] <= 8'h77;
		memory[16'h2233] <= 8'hd9;
		memory[16'h2234] <= 8'h46;
		memory[16'h2235] <= 8'h48;
		memory[16'h2236] <= 8'hec;
		memory[16'h2237] <= 8'h93;
		memory[16'h2238] <= 8'hb;
		memory[16'h2239] <= 8'hca;
		memory[16'h223a] <= 8'h44;
		memory[16'h223b] <= 8'h2a;
		memory[16'h223c] <= 8'hb1;
		memory[16'h223d] <= 8'hd3;
		memory[16'h223e] <= 8'h89;
		memory[16'h223f] <= 8'h20;
		memory[16'h2240] <= 8'h17;
		memory[16'h2241] <= 8'h21;
		memory[16'h2242] <= 8'hb2;
		memory[16'h2243] <= 8'had;
		memory[16'h2244] <= 8'h81;
		memory[16'h2245] <= 8'hd;
		memory[16'h2246] <= 8'h19;
		memory[16'h2247] <= 8'he6;
		memory[16'h2248] <= 8'h28;
		memory[16'h2249] <= 8'h77;
		memory[16'h224a] <= 8'haf;
		memory[16'h224b] <= 8'hbe;
		memory[16'h224c] <= 8'h1e;
		memory[16'h224d] <= 8'hd7;
		memory[16'h224e] <= 8'h2f;
		memory[16'h224f] <= 8'heb;
		memory[16'h2250] <= 8'hc;
		memory[16'h2251] <= 8'ha7;
		memory[16'h2252] <= 8'hc4;
		memory[16'h2253] <= 8'h53;
		memory[16'h2254] <= 8'hef;
		memory[16'h2255] <= 8'hb1;
		memory[16'h2256] <= 8'he6;
		memory[16'h2257] <= 8'hfa;
		memory[16'h2258] <= 8'h7b;
		memory[16'h2259] <= 8'h2a;
		memory[16'h225a] <= 8'h25;
		memory[16'h225b] <= 8'h2c;
		memory[16'h225c] <= 8'hfd;
		memory[16'h225d] <= 8'hae;
		memory[16'h225e] <= 8'h4d;
		memory[16'h225f] <= 8'h14;
		memory[16'h2260] <= 8'hcf;
		memory[16'h2261] <= 8'hff;
		memory[16'h2262] <= 8'hc2;
		memory[16'h2263] <= 8'h50;
		memory[16'h2264] <= 8'hc;
		memory[16'h2265] <= 8'hdb;
		memory[16'h2266] <= 8'h37;
		memory[16'h2267] <= 8'h34;
		memory[16'h2268] <= 8'h52;
		memory[16'h2269] <= 8'he6;
		memory[16'h226a] <= 8'hf2;
		memory[16'h226b] <= 8'h71;
		memory[16'h226c] <= 8'hbd;
		memory[16'h226d] <= 8'h21;
		memory[16'h226e] <= 8'h5c;
		memory[16'h226f] <= 8'hc9;
		memory[16'h2270] <= 8'hc8;
		memory[16'h2271] <= 8'h20;
		memory[16'h2272] <= 8'h1c;
		memory[16'h2273] <= 8'hb7;
		memory[16'h2274] <= 8'hd1;
		memory[16'h2275] <= 8'h2;
		memory[16'h2276] <= 8'hb2;
		memory[16'h2277] <= 8'h4d;
		memory[16'h2278] <= 8'h2c;
		memory[16'h2279] <= 8'hd7;
		memory[16'h227a] <= 8'h79;
		memory[16'h227b] <= 8'h29;
		memory[16'h227c] <= 8'h85;
		memory[16'h227d] <= 8'hc6;
		memory[16'h227e] <= 8'h3e;
		memory[16'h227f] <= 8'h55;
		memory[16'h2280] <= 8'hc5;
		memory[16'h2281] <= 8'h0;
		memory[16'h2282] <= 8'ha5;
		memory[16'h2283] <= 8'hd1;
		memory[16'h2284] <= 8'hdb;
		memory[16'h2285] <= 8'hdc;
		memory[16'h2286] <= 8'h5;
		memory[16'h2287] <= 8'h2e;
		memory[16'h2288] <= 8'hc2;
		memory[16'h2289] <= 8'hf7;
		memory[16'h228a] <= 8'h9f;
		memory[16'h228b] <= 8'h7f;
		memory[16'h228c] <= 8'h19;
		memory[16'h228d] <= 8'hfb;
		memory[16'h228e] <= 8'h49;
		memory[16'h228f] <= 8'he1;
		memory[16'h2290] <= 8'h1b;
		memory[16'h2291] <= 8'h65;
		memory[16'h2292] <= 8'h99;
		memory[16'h2293] <= 8'hed;
		memory[16'h2294] <= 8'h68;
		memory[16'h2295] <= 8'h4b;
		memory[16'h2296] <= 8'h3a;
		memory[16'h2297] <= 8'h94;
		memory[16'h2298] <= 8'h22;
		memory[16'h2299] <= 8'hb3;
		memory[16'h229a] <= 8'hbe;
		memory[16'h229b] <= 8'ha7;
		memory[16'h229c] <= 8'h7a;
		memory[16'h229d] <= 8'hfc;
		memory[16'h229e] <= 8'hfc;
		memory[16'h229f] <= 8'h3f;
		memory[16'h22a0] <= 8'hfc;
		memory[16'h22a1] <= 8'ha2;
		memory[16'h22a2] <= 8'h11;
		memory[16'h22a3] <= 8'hd7;
		memory[16'h22a4] <= 8'h7e;
		memory[16'h22a5] <= 8'h16;
		memory[16'h22a6] <= 8'h5;
		memory[16'h22a7] <= 8'h41;
		memory[16'h22a8] <= 8'he;
		memory[16'h22a9] <= 8'ha4;
		memory[16'h22aa] <= 8'hc0;
		memory[16'h22ab] <= 8'h27;
		memory[16'h22ac] <= 8'h9f;
		memory[16'h22ad] <= 8'h9;
		memory[16'h22ae] <= 8'h8;
		memory[16'h22af] <= 8'hbb;
		memory[16'h22b0] <= 8'h6f;
		memory[16'h22b1] <= 8'ha1;
		memory[16'h22b2] <= 8'ha8;
		memory[16'h22b3] <= 8'hd7;
		memory[16'h22b4] <= 8'hec;
		memory[16'h22b5] <= 8'he2;
		memory[16'h22b6] <= 8'h6b;
		memory[16'h22b7] <= 8'he;
		memory[16'h22b8] <= 8'h95;
		memory[16'h22b9] <= 8'h29;
		memory[16'h22ba] <= 8'hb6;
		memory[16'h22bb] <= 8'hf;
		memory[16'h22bc] <= 8'h25;
		memory[16'h22bd] <= 8'hb2;
		memory[16'h22be] <= 8'h4f;
		memory[16'h22bf] <= 8'h21;
		memory[16'h22c0] <= 8'h54;
		memory[16'h22c1] <= 8'h60;
		memory[16'h22c2] <= 8'hf9;
		memory[16'h22c3] <= 8'hd3;
		memory[16'h22c4] <= 8'h76;
		memory[16'h22c5] <= 8'hfe;
		memory[16'h22c6] <= 8'h14;
		memory[16'h22c7] <= 8'h84;
		memory[16'h22c8] <= 8'ha3;
		memory[16'h22c9] <= 8'hd4;
		memory[16'h22ca] <= 8'hab;
		memory[16'h22cb] <= 8'h42;
		memory[16'h22cc] <= 8'hde;
		memory[16'h22cd] <= 8'hb4;
		memory[16'h22ce] <= 8'hfd;
		memory[16'h22cf] <= 8'h4d;
		memory[16'h22d0] <= 8'h55;
		memory[16'h22d1] <= 8'ha5;
		memory[16'h22d2] <= 8'h24;
		memory[16'h22d3] <= 8'h42;
		memory[16'h22d4] <= 8'h87;
		memory[16'h22d5] <= 8'h8f;
		memory[16'h22d6] <= 8'h50;
		memory[16'h22d7] <= 8'h1d;
		memory[16'h22d8] <= 8'hb9;
		memory[16'h22d9] <= 8'h6;
		memory[16'h22da] <= 8'h2c;
		memory[16'h22db] <= 8'hde;
		memory[16'h22dc] <= 8'hb9;
		memory[16'h22dd] <= 8'h7b;
		memory[16'h22de] <= 8'h0;
		memory[16'h22df] <= 8'hd;
		memory[16'h22e0] <= 8'hdb;
		memory[16'h22e1] <= 8'hf9;
		memory[16'h22e2] <= 8'he0;
		memory[16'h22e3] <= 8'h52;
		memory[16'h22e4] <= 8'hf7;
		memory[16'h22e5] <= 8'hf4;
		memory[16'h22e6] <= 8'hd6;
		memory[16'h22e7] <= 8'h9a;
		memory[16'h22e8] <= 8'hc9;
		memory[16'h22e9] <= 8'h82;
		memory[16'h22ea] <= 8'hdd;
		memory[16'h22eb] <= 8'ha7;
		memory[16'h22ec] <= 8'h36;
		memory[16'h22ed] <= 8'hda;
		memory[16'h22ee] <= 8'hf4;
		memory[16'h22ef] <= 8'h8b;
		memory[16'h22f0] <= 8'h80;
		memory[16'h22f1] <= 8'h18;
		memory[16'h22f2] <= 8'hcd;
		memory[16'h22f3] <= 8'h7;
		memory[16'h22f4] <= 8'ha7;
		memory[16'h22f5] <= 8'h1e;
		memory[16'h22f6] <= 8'h24;
		memory[16'h22f7] <= 8'h60;
		memory[16'h22f8] <= 8'h24;
		memory[16'h22f9] <= 8'h51;
		memory[16'h22fa] <= 8'h3f;
		memory[16'h22fb] <= 8'hdd;
		memory[16'h22fc] <= 8'hcc;
		memory[16'h22fd] <= 8'h3f;
		memory[16'h22fe] <= 8'heb;
		memory[16'h22ff] <= 8'ha8;
		memory[16'h2300] <= 8'h38;
		memory[16'h2301] <= 8'hcb;
		memory[16'h2302] <= 8'hfa;
		memory[16'h2303] <= 8'h2f;
		memory[16'h2304] <= 8'hc0;
		memory[16'h2305] <= 8'hd0;
		memory[16'h2306] <= 8'hca;
		memory[16'h2307] <= 8'h89;
		memory[16'h2308] <= 8'h52;
		memory[16'h2309] <= 8'ha7;
		memory[16'h230a] <= 8'h30;
		memory[16'h230b] <= 8'h88;
		memory[16'h230c] <= 8'h81;
		memory[16'h230d] <= 8'h24;
		memory[16'h230e] <= 8'h14;
		memory[16'h230f] <= 8'h1;
		memory[16'h2310] <= 8'h3c;
		memory[16'h2311] <= 8'he1;
		memory[16'h2312] <= 8'h9;
		memory[16'h2313] <= 8'he3;
		memory[16'h2314] <= 8'hff;
		memory[16'h2315] <= 8'h2d;
		memory[16'h2316] <= 8'h44;
		memory[16'h2317] <= 8'h24;
		memory[16'h2318] <= 8'h7e;
		memory[16'h2319] <= 8'h83;
		memory[16'h231a] <= 8'h1;
		memory[16'h231b] <= 8'h4b;
		memory[16'h231c] <= 8'hc2;
		memory[16'h231d] <= 8'hec;
		memory[16'h231e] <= 8'hf3;
		memory[16'h231f] <= 8'hfa;
		memory[16'h2320] <= 8'hb8;
		memory[16'h2321] <= 8'hed;
		memory[16'h2322] <= 8'h29;
		memory[16'h2323] <= 8'h78;
		memory[16'h2324] <= 8'hbd;
		memory[16'h2325] <= 8'hf3;
		memory[16'h2326] <= 8'h1;
		memory[16'h2327] <= 8'h10;
		memory[16'h2328] <= 8'h9a;
		memory[16'h2329] <= 8'h31;
		memory[16'h232a] <= 8'h98;
		memory[16'h232b] <= 8'h1c;
		memory[16'h232c] <= 8'h55;
		memory[16'h232d] <= 8'hac;
		memory[16'h232e] <= 8'h1d;
		memory[16'h232f] <= 8'h91;
		memory[16'h2330] <= 8'h8e;
		memory[16'h2331] <= 8'h26;
		memory[16'h2332] <= 8'h74;
		memory[16'h2333] <= 8'h8d;
		memory[16'h2334] <= 8'h54;
		memory[16'h2335] <= 8'hb8;
		memory[16'h2336] <= 8'hb1;
		memory[16'h2337] <= 8'hd2;
		memory[16'h2338] <= 8'h3b;
		memory[16'h2339] <= 8'hb3;
		memory[16'h233a] <= 8'h1d;
		memory[16'h233b] <= 8'hfd;
		memory[16'h233c] <= 8'h9f;
		memory[16'h233d] <= 8'h10;
		memory[16'h233e] <= 8'hf7;
		memory[16'h233f] <= 8'h57;
		memory[16'h2340] <= 8'hfd;
		memory[16'h2341] <= 8'h21;
		memory[16'h2342] <= 8'hcf;
		memory[16'h2343] <= 8'hbb;
		memory[16'h2344] <= 8'h14;
		memory[16'h2345] <= 8'hd0;
		memory[16'h2346] <= 8'hcb;
		memory[16'h2347] <= 8'haf;
		memory[16'h2348] <= 8'h1;
		memory[16'h2349] <= 8'h63;
		memory[16'h234a] <= 8'hcb;
		memory[16'h234b] <= 8'h56;
		memory[16'h234c] <= 8'h10;
		memory[16'h234d] <= 8'he8;
		memory[16'h234e] <= 8'he7;
		memory[16'h234f] <= 8'h9e;
		memory[16'h2350] <= 8'hf;
		memory[16'h2351] <= 8'h5c;
		memory[16'h2352] <= 8'h2b;
		memory[16'h2353] <= 8'h63;
		memory[16'h2354] <= 8'h14;
		memory[16'h2355] <= 8'hdd;
		memory[16'h2356] <= 8'h35;
		memory[16'h2357] <= 8'h50;
		memory[16'h2358] <= 8'h90;
		memory[16'h2359] <= 8'h53;
		memory[16'h235a] <= 8'h4d;
		memory[16'h235b] <= 8'h2f;
		memory[16'h235c] <= 8'h63;
		memory[16'h235d] <= 8'h45;
		memory[16'h235e] <= 8'h87;
		memory[16'h235f] <= 8'h61;
		memory[16'h2360] <= 8'h66;
		memory[16'h2361] <= 8'h56;
		memory[16'h2362] <= 8'h1c;
		memory[16'h2363] <= 8'h7a;
		memory[16'h2364] <= 8'h27;
		memory[16'h2365] <= 8'he7;
		memory[16'h2366] <= 8'h29;
		memory[16'h2367] <= 8'h28;
		memory[16'h2368] <= 8'h4a;
		memory[16'h2369] <= 8'hf4;
		memory[16'h236a] <= 8'h7f;
		memory[16'h236b] <= 8'h5a;
		memory[16'h236c] <= 8'hdd;
		memory[16'h236d] <= 8'h66;
		memory[16'h236e] <= 8'hf8;
		memory[16'h236f] <= 8'hec;
		memory[16'h2370] <= 8'hc2;
		memory[16'h2371] <= 8'h24;
		memory[16'h2372] <= 8'h4f;
		memory[16'h2373] <= 8'hd7;
		memory[16'h2374] <= 8'h1;
		memory[16'h2375] <= 8'h84;
		memory[16'h2376] <= 8'h27;
		memory[16'h2377] <= 8'h91;
		memory[16'h2378] <= 8'hd7;
		memory[16'h2379] <= 8'h74;
		memory[16'h237a] <= 8'hc0;
		memory[16'h237b] <= 8'h3b;
		memory[16'h237c] <= 8'hb9;
		memory[16'h237d] <= 8'h47;
		memory[16'h237e] <= 8'h9c;
		memory[16'h237f] <= 8'h1f;
		memory[16'h2380] <= 8'h9e;
		memory[16'h2381] <= 8'hb8;
		memory[16'h2382] <= 8'h9a;
		memory[16'h2383] <= 8'hc5;
		memory[16'h2384] <= 8'h9f;
		memory[16'h2385] <= 8'hc3;
		memory[16'h2386] <= 8'hed;
		memory[16'h2387] <= 8'he9;
		memory[16'h2388] <= 8'hb8;
		memory[16'h2389] <= 8'h6c;
		memory[16'h238a] <= 8'h44;
		memory[16'h238b] <= 8'h95;
		memory[16'h238c] <= 8'hd3;
		memory[16'h238d] <= 8'h3c;
		memory[16'h238e] <= 8'h81;
		memory[16'h238f] <= 8'h95;
		memory[16'h2390] <= 8'h60;
		memory[16'h2391] <= 8'hd0;
		memory[16'h2392] <= 8'h6c;
		memory[16'h2393] <= 8'h61;
		memory[16'h2394] <= 8'h54;
		memory[16'h2395] <= 8'h93;
		memory[16'h2396] <= 8'hf2;
		memory[16'h2397] <= 8'h2c;
		memory[16'h2398] <= 8'h8;
		memory[16'h2399] <= 8'hb3;
		memory[16'h239a] <= 8'h67;
		memory[16'h239b] <= 8'hc1;
		memory[16'h239c] <= 8'hfa;
		memory[16'h239d] <= 8'h3;
		memory[16'h239e] <= 8'he1;
		memory[16'h239f] <= 8'h98;
		memory[16'h23a0] <= 8'hbb;
		memory[16'h23a1] <= 8'h7b;
		memory[16'h23a2] <= 8'h5d;
		memory[16'h23a3] <= 8'h5a;
		memory[16'h23a4] <= 8'h3e;
		memory[16'h23a5] <= 8'h4b;
		memory[16'h23a6] <= 8'h43;
		memory[16'h23a7] <= 8'hf6;
		memory[16'h23a8] <= 8'hb7;
		memory[16'h23a9] <= 8'h87;
		memory[16'h23aa] <= 8'h8b;
		memory[16'h23ab] <= 8'h8a;
		memory[16'h23ac] <= 8'hc4;
		memory[16'h23ad] <= 8'hc;
		memory[16'h23ae] <= 8'h20;
		memory[16'h23af] <= 8'h24;
		memory[16'h23b0] <= 8'hdc;
		memory[16'h23b1] <= 8'h8c;
		memory[16'h23b2] <= 8'h86;
		memory[16'h23b3] <= 8'h31;
		memory[16'h23b4] <= 8'h20;
		memory[16'h23b5] <= 8'h78;
		memory[16'h23b6] <= 8'h5d;
		memory[16'h23b7] <= 8'h28;
		memory[16'h23b8] <= 8'h2b;
		memory[16'h23b9] <= 8'hc4;
		memory[16'h23ba] <= 8'he9;
		memory[16'h23bb] <= 8'h26;
		memory[16'h23bc] <= 8'hc7;
		memory[16'h23bd] <= 8'hca;
		memory[16'h23be] <= 8'hbe;
		memory[16'h23bf] <= 8'h82;
		memory[16'h23c0] <= 8'h45;
		memory[16'h23c1] <= 8'h1c;
		memory[16'h23c2] <= 8'hdc;
		memory[16'h23c3] <= 8'h84;
		memory[16'h23c4] <= 8'h67;
		memory[16'h23c5] <= 8'h1f;
		memory[16'h23c6] <= 8'h7a;
		memory[16'h23c7] <= 8'h1e;
		memory[16'h23c8] <= 8'ha7;
		memory[16'h23c9] <= 8'h6;
		memory[16'h23ca] <= 8'ha9;
		memory[16'h23cb] <= 8'h6b;
		memory[16'h23cc] <= 8'h12;
		memory[16'h23cd] <= 8'hc9;
		memory[16'h23ce] <= 8'h8f;
		memory[16'h23cf] <= 8'hef;
		memory[16'h23d0] <= 8'h55;
		memory[16'h23d1] <= 8'h15;
		memory[16'h23d2] <= 8'h20;
		memory[16'h23d3] <= 8'h75;
		memory[16'h23d4] <= 8'h8e;
		memory[16'h23d5] <= 8'h7d;
		memory[16'h23d6] <= 8'h9d;
		memory[16'h23d7] <= 8'hb9;
		memory[16'h23d8] <= 8'h41;
		memory[16'h23d9] <= 8'h87;
		memory[16'h23da] <= 8'hdf;
		memory[16'h23db] <= 8'h8;
		memory[16'h23dc] <= 8'h51;
		memory[16'h23dd] <= 8'h9e;
		memory[16'h23de] <= 8'h8a;
		memory[16'h23df] <= 8'h97;
		memory[16'h23e0] <= 8'hba;
		memory[16'h23e1] <= 8'h66;
		memory[16'h23e2] <= 8'h1b;
		memory[16'h23e3] <= 8'h21;
		memory[16'h23e4] <= 8'h85;
		memory[16'h23e5] <= 8'h95;
		memory[16'h23e6] <= 8'h3f;
		memory[16'h23e7] <= 8'h2c;
		memory[16'h23e8] <= 8'h9b;
		memory[16'h23e9] <= 8'he8;
		memory[16'h23ea] <= 8'h97;
		memory[16'h23eb] <= 8'hae;
		memory[16'h23ec] <= 8'hb1;
		memory[16'h23ed] <= 8'h27;
		memory[16'h23ee] <= 8'h9d;
		memory[16'h23ef] <= 8'h7;
		memory[16'h23f0] <= 8'h3c;
		memory[16'h23f1] <= 8'hbd;
		memory[16'h23f2] <= 8'h7c;
		memory[16'h23f3] <= 8'hca;
		memory[16'h23f4] <= 8'h3a;
		memory[16'h23f5] <= 8'h1a;
		memory[16'h23f6] <= 8'h84;
		memory[16'h23f7] <= 8'h7b;
		memory[16'h23f8] <= 8'ha1;
		memory[16'h23f9] <= 8'h63;
		memory[16'h23fa] <= 8'h83;
		memory[16'h23fb] <= 8'hf2;
		memory[16'h23fc] <= 8'h1;
		memory[16'h23fd] <= 8'hd;
		memory[16'h23fe] <= 8'h89;
		memory[16'h23ff] <= 8'hbb;
		memory[16'h2400] <= 8'h73;
		memory[16'h2401] <= 8'ha4;
		memory[16'h2402] <= 8'hdc;
		memory[16'h2403] <= 8'hf8;
		memory[16'h2404] <= 8'h3a;
		memory[16'h2405] <= 8'h1c;
		memory[16'h2406] <= 8'h25;
		memory[16'h2407] <= 8'hd5;
		memory[16'h2408] <= 8'h4;
		memory[16'h2409] <= 8'hbc;
		memory[16'h240a] <= 8'h83;
		memory[16'h240b] <= 8'hb6;
		memory[16'h240c] <= 8'he3;
		memory[16'h240d] <= 8'h20;
		memory[16'h240e] <= 8'hbd;
		memory[16'h240f] <= 8'h20;
		memory[16'h2410] <= 8'hdd;
		memory[16'h2411] <= 8'h39;
		memory[16'h2412] <= 8'hea;
		memory[16'h2413] <= 8'h17;
		memory[16'h2414] <= 8'h53;
		memory[16'h2415] <= 8'h6e;
		memory[16'h2416] <= 8'h92;
		memory[16'h2417] <= 8'hf4;
		memory[16'h2418] <= 8'hd2;
		memory[16'h2419] <= 8'h15;
		memory[16'h241a] <= 8'he7;
		memory[16'h241b] <= 8'hd3;
		memory[16'h241c] <= 8'h22;
		memory[16'h241d] <= 8'h70;
		memory[16'h241e] <= 8'h8f;
		memory[16'h241f] <= 8'h95;
		memory[16'h2420] <= 8'h15;
		memory[16'h2421] <= 8'h6b;
		memory[16'h2422] <= 8'h8e;
		memory[16'h2423] <= 8'h4f;
		memory[16'h2424] <= 8'h87;
		memory[16'h2425] <= 8'hb3;
		memory[16'h2426] <= 8'h24;
		memory[16'h2427] <= 8'h8c;
		memory[16'h2428] <= 8'h6f;
		memory[16'h2429] <= 8'ha8;
		memory[16'h242a] <= 8'h42;
		memory[16'h242b] <= 8'h53;
		memory[16'h242c] <= 8'hc8;
		memory[16'h242d] <= 8'hff;
		memory[16'h242e] <= 8'h73;
		memory[16'h242f] <= 8'ha6;
		memory[16'h2430] <= 8'h38;
		memory[16'h2431] <= 8'h5d;
		memory[16'h2432] <= 8'hbd;
		memory[16'h2433] <= 8'h8c;
		memory[16'h2434] <= 8'hcc;
		memory[16'h2435] <= 8'h50;
		memory[16'h2436] <= 8'h80;
		memory[16'h2437] <= 8'h9e;
		memory[16'h2438] <= 8'h65;
		memory[16'h2439] <= 8'h67;
		memory[16'h243a] <= 8'h71;
		memory[16'h243b] <= 8'h88;
		memory[16'h243c] <= 8'hd8;
		memory[16'h243d] <= 8'h0;
		memory[16'h243e] <= 8'h1d;
		memory[16'h243f] <= 8'hed;
		memory[16'h2440] <= 8'h6c;
		memory[16'h2441] <= 8'hab;
		memory[16'h2442] <= 8'h3c;
		memory[16'h2443] <= 8'hf3;
		memory[16'h2444] <= 8'h5e;
		memory[16'h2445] <= 8'h60;
		memory[16'h2446] <= 8'h7f;
		memory[16'h2447] <= 8'hce;
		memory[16'h2448] <= 8'h8;
		memory[16'h2449] <= 8'hc1;
		memory[16'h244a] <= 8'h21;
		memory[16'h244b] <= 8'hd1;
		memory[16'h244c] <= 8'hc0;
		memory[16'h244d] <= 8'h94;
		memory[16'h244e] <= 8'h77;
		memory[16'h244f] <= 8'hf9;
		memory[16'h2450] <= 8'hf1;
		memory[16'h2451] <= 8'h34;
		memory[16'h2452] <= 8'h85;
		memory[16'h2453] <= 8'hbd;
		memory[16'h2454] <= 8'h84;
		memory[16'h2455] <= 8'h5;
		memory[16'h2456] <= 8'h5b;
		memory[16'h2457] <= 8'hea;
		memory[16'h2458] <= 8'h6d;
		memory[16'h2459] <= 8'hcd;
		memory[16'h245a] <= 8'h72;
		memory[16'h245b] <= 8'h45;
		memory[16'h245c] <= 8'hcd;
		memory[16'h245d] <= 8'h8f;
		memory[16'h245e] <= 8'h32;
		memory[16'h245f] <= 8'h39;
		memory[16'h2460] <= 8'h3b;
		memory[16'h2461] <= 8'h6e;
		memory[16'h2462] <= 8'h2d;
		memory[16'h2463] <= 8'h99;
		memory[16'h2464] <= 8'hce;
		memory[16'h2465] <= 8'hac;
		memory[16'h2466] <= 8'h67;
		memory[16'h2467] <= 8'hd7;
		memory[16'h2468] <= 8'h6e;
		memory[16'h2469] <= 8'h88;
		memory[16'h246a] <= 8'ha8;
		memory[16'h246b] <= 8'h2e;
		memory[16'h246c] <= 8'h1c;
		memory[16'h246d] <= 8'h1f;
		memory[16'h246e] <= 8'h27;
		memory[16'h246f] <= 8'he;
		memory[16'h2470] <= 8'h53;
		memory[16'h2471] <= 8'hac;
		memory[16'h2472] <= 8'hcb;
		memory[16'h2473] <= 8'hd8;
		memory[16'h2474] <= 8'hb2;
		memory[16'h2475] <= 8'h27;
		memory[16'h2476] <= 8'hc2;
		memory[16'h2477] <= 8'h1f;
		memory[16'h2478] <= 8'hf4;
		memory[16'h2479] <= 8'h34;
		memory[16'h247a] <= 8'h64;
		memory[16'h247b] <= 8'hc1;
		memory[16'h247c] <= 8'hc3;
		memory[16'h247d] <= 8'h96;
		memory[16'h247e] <= 8'hfb;
		memory[16'h247f] <= 8'hfe;
		memory[16'h2480] <= 8'h4;
		memory[16'h2481] <= 8'h28;
		memory[16'h2482] <= 8'h98;
		memory[16'h2483] <= 8'hd2;
		memory[16'h2484] <= 8'hd4;
		memory[16'h2485] <= 8'hff;
		memory[16'h2486] <= 8'ha9;
		memory[16'h2487] <= 8'h42;
		memory[16'h2488] <= 8'h88;
		memory[16'h2489] <= 8'h51;
		memory[16'h248a] <= 8'h71;
		memory[16'h248b] <= 8'ha4;
		memory[16'h248c] <= 8'h70;
		memory[16'h248d] <= 8'h98;
		memory[16'h248e] <= 8'hb2;
		memory[16'h248f] <= 8'hc4;
		memory[16'h2490] <= 8'h45;
		memory[16'h2491] <= 8'h7e;
		memory[16'h2492] <= 8'h9c;
		memory[16'h2493] <= 8'hf7;
		memory[16'h2494] <= 8'ha5;
		memory[16'h2495] <= 8'h5e;
		memory[16'h2496] <= 8'h16;
		memory[16'h2497] <= 8'h99;
		memory[16'h2498] <= 8'h92;
		memory[16'h2499] <= 8'h7a;
		memory[16'h249a] <= 8'h5a;
		memory[16'h249b] <= 8'h55;
		memory[16'h249c] <= 8'h10;
		memory[16'h249d] <= 8'h55;
		memory[16'h249e] <= 8'h54;
		memory[16'h249f] <= 8'h14;
		memory[16'h24a0] <= 8'h7d;
		memory[16'h24a1] <= 8'hec;
		memory[16'h24a2] <= 8'he6;
		memory[16'h24a3] <= 8'h52;
		memory[16'h24a4] <= 8'heb;
		memory[16'h24a5] <= 8'h90;
		memory[16'h24a6] <= 8'h94;
		memory[16'h24a7] <= 8'h73;
		memory[16'h24a8] <= 8'he1;
		memory[16'h24a9] <= 8'h5;
		memory[16'h24aa] <= 8'h18;
		memory[16'h24ab] <= 8'h52;
		memory[16'h24ac] <= 8'h9e;
		memory[16'h24ad] <= 8'hca;
		memory[16'h24ae] <= 8'h16;
		memory[16'h24af] <= 8'he3;
		memory[16'h24b0] <= 8'h48;
		memory[16'h24b1] <= 8'hb2;
		memory[16'h24b2] <= 8'hda;
		memory[16'h24b3] <= 8'hed;
		memory[16'h24b4] <= 8'h10;
		memory[16'h24b5] <= 8'hf0;
		memory[16'h24b6] <= 8'h86;
		memory[16'h24b7] <= 8'ha2;
		memory[16'h24b8] <= 8'h6a;
		memory[16'h24b9] <= 8'he1;
		memory[16'h24ba] <= 8'hf7;
		memory[16'h24bb] <= 8'h7a;
		memory[16'h24bc] <= 8'h36;
		memory[16'h24bd] <= 8'h4b;
		memory[16'h24be] <= 8'h8e;
		memory[16'h24bf] <= 8'hb4;
		memory[16'h24c0] <= 8'h37;
		memory[16'h24c1] <= 8'h74;
		memory[16'h24c2] <= 8'h6;
		memory[16'h24c3] <= 8'h23;
		memory[16'h24c4] <= 8'h4;
		memory[16'h24c5] <= 8'h9a;
		memory[16'h24c6] <= 8'h96;
		memory[16'h24c7] <= 8'he6;
		memory[16'h24c8] <= 8'ha0;
		memory[16'h24c9] <= 8'hae;
		memory[16'h24ca] <= 8'h38;
		memory[16'h24cb] <= 8'h3e;
		memory[16'h24cc] <= 8'h79;
		memory[16'h24cd] <= 8'h4e;
		memory[16'h24ce] <= 8'h21;
		memory[16'h24cf] <= 8'hc1;
		memory[16'h24d0] <= 8'h0;
		memory[16'h24d1] <= 8'hfb;
		memory[16'h24d2] <= 8'haf;
		memory[16'h24d3] <= 8'h10;
		memory[16'h24d4] <= 8'heb;
		memory[16'h24d5] <= 8'h35;
		memory[16'h24d6] <= 8'hb2;
		memory[16'h24d7] <= 8'h55;
		memory[16'h24d8] <= 8'h16;
		memory[16'h24d9] <= 8'ha9;
		memory[16'h24da] <= 8'hcf;
		memory[16'h24db] <= 8'h4d;
		memory[16'h24dc] <= 8'hf5;
		memory[16'h24dd] <= 8'h5d;
		memory[16'h24de] <= 8'h1;
		memory[16'h24df] <= 8'h2c;
		memory[16'h24e0] <= 8'hd1;
		memory[16'h24e1] <= 8'h7;
		memory[16'h24e2] <= 8'h4f;
		memory[16'h24e3] <= 8'hd6;
		memory[16'h24e4] <= 8'ha1;
		memory[16'h24e5] <= 8'he6;
		memory[16'h24e6] <= 8'hbc;
		memory[16'h24e7] <= 8'h41;
		memory[16'h24e8] <= 8'h94;
		memory[16'h24e9] <= 8'hf4;
		memory[16'h24ea] <= 8'h7f;
		memory[16'h24eb] <= 8'hd;
		memory[16'h24ec] <= 8'h42;
		memory[16'h24ed] <= 8'ha0;
		memory[16'h24ee] <= 8'hcf;
		memory[16'h24ef] <= 8'h42;
		memory[16'h24f0] <= 8'h9b;
		memory[16'h24f1] <= 8'h7e;
		memory[16'h24f2] <= 8'h52;
		memory[16'h24f3] <= 8'h86;
		memory[16'h24f4] <= 8'hb3;
		memory[16'h24f5] <= 8'h4;
		memory[16'h24f6] <= 8'hdb;
		memory[16'h24f7] <= 8'hca;
		memory[16'h24f8] <= 8'had;
		memory[16'h24f9] <= 8'haa;
		memory[16'h24fa] <= 8'h17;
		memory[16'h24fb] <= 8'ha2;
		memory[16'h24fc] <= 8'h7;
		memory[16'h24fd] <= 8'h18;
		memory[16'h24fe] <= 8'hcf;
		memory[16'h24ff] <= 8'hd9;
		memory[16'h2500] <= 8'h1f;
		memory[16'h2501] <= 8'h1e;
		memory[16'h2502] <= 8'haf;
		memory[16'h2503] <= 8'hc0;
		memory[16'h2504] <= 8'h4;
		memory[16'h2505] <= 8'h6b;
		memory[16'h2506] <= 8'h2;
		memory[16'h2507] <= 8'h99;
		memory[16'h2508] <= 8'h5f;
		memory[16'h2509] <= 8'h81;
		memory[16'h250a] <= 8'ha6;
		memory[16'h250b] <= 8'ha1;
		memory[16'h250c] <= 8'h22;
		memory[16'h250d] <= 8'h75;
		memory[16'h250e] <= 8'he3;
		memory[16'h250f] <= 8'hbd;
		memory[16'h2510] <= 8'hf3;
		memory[16'h2511] <= 8'h35;
		memory[16'h2512] <= 8'h44;
		memory[16'h2513] <= 8'ha7;
		memory[16'h2514] <= 8'h39;
		memory[16'h2515] <= 8'h1f;
		memory[16'h2516] <= 8'h71;
		memory[16'h2517] <= 8'he6;
		memory[16'h2518] <= 8'hca;
		memory[16'h2519] <= 8'h88;
		memory[16'h251a] <= 8'h89;
		memory[16'h251b] <= 8'hd1;
		memory[16'h251c] <= 8'ha0;
		memory[16'h251d] <= 8'h58;
		memory[16'h251e] <= 8'haa;
		memory[16'h251f] <= 8'hbf;
		memory[16'h2520] <= 8'h76;
		memory[16'h2521] <= 8'h59;
		memory[16'h2522] <= 8'h7f;
		memory[16'h2523] <= 8'h7b;
		memory[16'h2524] <= 8'hc4;
		memory[16'h2525] <= 8'h81;
		memory[16'h2526] <= 8'h14;
		memory[16'h2527] <= 8'h23;
		memory[16'h2528] <= 8'h3;
		memory[16'h2529] <= 8'hba;
		memory[16'h252a] <= 8'hc4;
		memory[16'h252b] <= 8'h25;
		memory[16'h252c] <= 8'h30;
		memory[16'h252d] <= 8'ha7;
		memory[16'h252e] <= 8'he2;
		memory[16'h252f] <= 8'h23;
		memory[16'h2530] <= 8'hdc;
		memory[16'h2531] <= 8'h26;
		memory[16'h2532] <= 8'hca;
		memory[16'h2533] <= 8'h15;
		memory[16'h2534] <= 8'h46;
		memory[16'h2535] <= 8'h3b;
		memory[16'h2536] <= 8'hfc;
		memory[16'h2537] <= 8'h10;
		memory[16'h2538] <= 8'hc3;
		memory[16'h2539] <= 8'h85;
		memory[16'h253a] <= 8'he1;
		memory[16'h253b] <= 8'h63;
		memory[16'h253c] <= 8'hdd;
		memory[16'h253d] <= 8'h8c;
		memory[16'h253e] <= 8'h22;
		memory[16'h253f] <= 8'h53;
		memory[16'h2540] <= 8'he5;
		memory[16'h2541] <= 8'ha2;
		memory[16'h2542] <= 8'hce;
		memory[16'h2543] <= 8'haa;
		memory[16'h2544] <= 8'h23;
		memory[16'h2545] <= 8'he2;
		memory[16'h2546] <= 8'hcd;
		memory[16'h2547] <= 8'h26;
		memory[16'h2548] <= 8'h9d;
		memory[16'h2549] <= 8'h92;
		memory[16'h254a] <= 8'h4b;
		memory[16'h254b] <= 8'hcd;
		memory[16'h254c] <= 8'h39;
		memory[16'h254d] <= 8'h2e;
		memory[16'h254e] <= 8'hf0;
		memory[16'h254f] <= 8'h16;
		memory[16'h2550] <= 8'h54;
		memory[16'h2551] <= 8'hbb;
		memory[16'h2552] <= 8'h2b;
		memory[16'h2553] <= 8'h9a;
		memory[16'h2554] <= 8'hf6;
		memory[16'h2555] <= 8'h27;
		memory[16'h2556] <= 8'haa;
		memory[16'h2557] <= 8'hba;
		memory[16'h2558] <= 8'hac;
		memory[16'h2559] <= 8'h8c;
		memory[16'h255a] <= 8'h1d;
		memory[16'h255b] <= 8'h89;
		memory[16'h255c] <= 8'h18;
		memory[16'h255d] <= 8'h40;
		memory[16'h255e] <= 8'hdd;
		memory[16'h255f] <= 8'hfd;
		memory[16'h2560] <= 8'he2;
		memory[16'h2561] <= 8'hab;
		memory[16'h2562] <= 8'ha7;
		memory[16'h2563] <= 8'h5;
		memory[16'h2564] <= 8'h8e;
		memory[16'h2565] <= 8'h75;
		memory[16'h2566] <= 8'h2c;
		memory[16'h2567] <= 8'h2b;
		memory[16'h2568] <= 8'h7;
		memory[16'h2569] <= 8'h77;
		memory[16'h256a] <= 8'hf8;
		memory[16'h256b] <= 8'h40;
		memory[16'h256c] <= 8'ha5;
		memory[16'h256d] <= 8'he8;
		memory[16'h256e] <= 8'h56;
		memory[16'h256f] <= 8'hfa;
		memory[16'h2570] <= 8'ha3;
		memory[16'h2571] <= 8'h82;
		memory[16'h2572] <= 8'h94;
		memory[16'h2573] <= 8'h9a;
		memory[16'h2574] <= 8'ha9;
		memory[16'h2575] <= 8'h3f;
		memory[16'h2576] <= 8'h54;
		memory[16'h2577] <= 8'h56;
		memory[16'h2578] <= 8'hcb;
		memory[16'h2579] <= 8'h71;
		memory[16'h257a] <= 8'hdf;
		memory[16'h257b] <= 8'he3;
		memory[16'h257c] <= 8'hb1;
		memory[16'h257d] <= 8'hbc;
		memory[16'h257e] <= 8'he0;
		memory[16'h257f] <= 8'h93;
		memory[16'h2580] <= 8'h68;
		memory[16'h2581] <= 8'h88;
		memory[16'h2582] <= 8'h99;
		memory[16'h2583] <= 8'hf6;
		memory[16'h2584] <= 8'hfd;
		memory[16'h2585] <= 8'hc5;
		memory[16'h2586] <= 8'h21;
		memory[16'h2587] <= 8'h4;
		memory[16'h2588] <= 8'h3c;
		memory[16'h2589] <= 8'h19;
		memory[16'h258a] <= 8'h44;
		memory[16'h258b] <= 8'he2;
		memory[16'h258c] <= 8'h1;
		memory[16'h258d] <= 8'h9b;
		memory[16'h258e] <= 8'hdc;
		memory[16'h258f] <= 8'ha5;
		memory[16'h2590] <= 8'h1d;
		memory[16'h2591] <= 8'h70;
		memory[16'h2592] <= 8'h3f;
		memory[16'h2593] <= 8'hc6;
		memory[16'h2594] <= 8'haf;
		memory[16'h2595] <= 8'h93;
		memory[16'h2596] <= 8'h1c;
		memory[16'h2597] <= 8'h7a;
		memory[16'h2598] <= 8'h4;
		memory[16'h2599] <= 8'hfc;
		memory[16'h259a] <= 8'h5d;
		memory[16'h259b] <= 8'hb6;
		memory[16'h259c] <= 8'hb8;
		memory[16'h259d] <= 8'h3e;
		memory[16'h259e] <= 8'h49;
		memory[16'h259f] <= 8'h20;
		memory[16'h25a0] <= 8'hc6;
		memory[16'h25a1] <= 8'he2;
		memory[16'h25a2] <= 8'h16;
		memory[16'h25a3] <= 8'hc3;
		memory[16'h25a4] <= 8'ha7;
		memory[16'h25a5] <= 8'h37;
		memory[16'h25a6] <= 8'hc7;
		memory[16'h25a7] <= 8'he4;
		memory[16'h25a8] <= 8'h50;
		memory[16'h25a9] <= 8'hb;
		memory[16'h25aa] <= 8'hc6;
		memory[16'h25ab] <= 8'h52;
		memory[16'h25ac] <= 8'ha6;
		memory[16'h25ad] <= 8'ha2;
		memory[16'h25ae] <= 8'hf7;
		memory[16'h25af] <= 8'hc3;
		memory[16'h25b0] <= 8'h12;
		memory[16'h25b1] <= 8'h36;
		memory[16'h25b2] <= 8'h8a;
		memory[16'h25b3] <= 8'hc2;
		memory[16'h25b4] <= 8'hc9;
		memory[16'h25b5] <= 8'ha6;
		memory[16'h25b6] <= 8'h3c;
		memory[16'h25b7] <= 8'hcd;
		memory[16'h25b8] <= 8'ha2;
		memory[16'h25b9] <= 8'h9a;
		memory[16'h25ba] <= 8'h83;
		memory[16'h25bb] <= 8'h5b;
		memory[16'h25bc] <= 8'hd8;
		memory[16'h25bd] <= 8'hcd;
		memory[16'h25be] <= 8'h7b;
		memory[16'h25bf] <= 8'h9e;
		memory[16'h25c0] <= 8'haf;
		memory[16'h25c1] <= 8'h92;
		memory[16'h25c2] <= 8'h61;
		memory[16'h25c3] <= 8'h57;
		memory[16'h25c4] <= 8'hc9;
		memory[16'h25c5] <= 8'h28;
		memory[16'h25c6] <= 8'h3b;
		memory[16'h25c7] <= 8'h1a;
		memory[16'h25c8] <= 8'h33;
		memory[16'h25c9] <= 8'h1;
		memory[16'h25ca] <= 8'h6c;
		memory[16'h25cb] <= 8'hda;
		memory[16'h25cc] <= 8'ha3;
		memory[16'h25cd] <= 8'h63;
		memory[16'h25ce] <= 8'h9d;
		memory[16'h25cf] <= 8'hb5;
		memory[16'h25d0] <= 8'h99;
		memory[16'h25d1] <= 8'h27;
		memory[16'h25d2] <= 8'h77;
		memory[16'h25d3] <= 8'h62;
		memory[16'h25d4] <= 8'hce;
		memory[16'h25d5] <= 8'hb4;
		memory[16'h25d6] <= 8'h2f;
		memory[16'h25d7] <= 8'h70;
		memory[16'h25d8] <= 8'h4e;
		memory[16'h25d9] <= 8'hb3;
		memory[16'h25da] <= 8'hcb;
		memory[16'h25db] <= 8'h26;
		memory[16'h25dc] <= 8'h80;
		memory[16'h25dd] <= 8'h47;
		memory[16'h25de] <= 8'hc4;
		memory[16'h25df] <= 8'h2f;
		memory[16'h25e0] <= 8'hd9;
		memory[16'h25e1] <= 8'h25;
		memory[16'h25e2] <= 8'h86;
		memory[16'h25e3] <= 8'ha2;
		memory[16'h25e4] <= 8'h4d;
		memory[16'h25e5] <= 8'hc1;
		memory[16'h25e6] <= 8'hbc;
		memory[16'h25e7] <= 8'h80;
		memory[16'h25e8] <= 8'hc2;
		memory[16'h25e9] <= 8'h28;
		memory[16'h25ea] <= 8'h5a;
		memory[16'h25eb] <= 8'h65;
		memory[16'h25ec] <= 8'h8b;
		memory[16'h25ed] <= 8'hf8;
		memory[16'h25ee] <= 8'h1b;
		memory[16'h25ef] <= 8'h24;
		memory[16'h25f0] <= 8'h1f;
		memory[16'h25f1] <= 8'h92;
		memory[16'h25f2] <= 8'h86;
		memory[16'h25f3] <= 8'hed;
		memory[16'h25f4] <= 8'h46;
		memory[16'h25f5] <= 8'hb6;
		memory[16'h25f6] <= 8'h5e;
		memory[16'h25f7] <= 8'h94;
		memory[16'h25f8] <= 8'h69;
		memory[16'h25f9] <= 8'h29;
		memory[16'h25fa] <= 8'hba;
		memory[16'h25fb] <= 8'he9;
		memory[16'h25fc] <= 8'h70;
		memory[16'h25fd] <= 8'h7e;
		memory[16'h25fe] <= 8'h18;
		memory[16'h25ff] <= 8'h49;
		memory[16'h2600] <= 8'ha3;
		memory[16'h2601] <= 8'h9f;
		memory[16'h2602] <= 8'hec;
		memory[16'h2603] <= 8'hf0;
		memory[16'h2604] <= 8'h60;
		memory[16'h2605] <= 8'ha8;
		memory[16'h2606] <= 8'h71;
		memory[16'h2607] <= 8'h23;
		memory[16'h2608] <= 8'hd1;
		memory[16'h2609] <= 8'hcb;
		memory[16'h260a] <= 8'h88;
		memory[16'h260b] <= 8'h5c;
		memory[16'h260c] <= 8'hc3;
		memory[16'h260d] <= 8'ha3;
		memory[16'h260e] <= 8'h81;
		memory[16'h260f] <= 8'he3;
		memory[16'h2610] <= 8'h36;
		memory[16'h2611] <= 8'h7;
		memory[16'h2612] <= 8'hd0;
		memory[16'h2613] <= 8'h7c;
		memory[16'h2614] <= 8'hbd;
		memory[16'h2615] <= 8'h2e;
		memory[16'h2616] <= 8'h11;
		memory[16'h2617] <= 8'h26;
		memory[16'h2618] <= 8'h58;
		memory[16'h2619] <= 8'hcb;
		memory[16'h261a] <= 8'hf;
		memory[16'h261b] <= 8'hc8;
		memory[16'h261c] <= 8'h4a;
		memory[16'h261d] <= 8'h28;
		memory[16'h261e] <= 8'h12;
		memory[16'h261f] <= 8'hed;
		memory[16'h2620] <= 8'hc7;
		memory[16'h2621] <= 8'hfe;
		memory[16'h2622] <= 8'hde;
		memory[16'h2623] <= 8'h27;
		memory[16'h2624] <= 8'ha6;
		memory[16'h2625] <= 8'h4f;
		memory[16'h2626] <= 8'h4a;
		memory[16'h2627] <= 8'h77;
		memory[16'h2628] <= 8'h1a;
		memory[16'h2629] <= 8'hd3;
		memory[16'h262a] <= 8'hd4;
		memory[16'h262b] <= 8'hde;
		memory[16'h262c] <= 8'h76;
		memory[16'h262d] <= 8'h55;
		memory[16'h262e] <= 8'hc1;
		memory[16'h262f] <= 8'hac;
		memory[16'h2630] <= 8'h5c;
		memory[16'h2631] <= 8'h91;
		memory[16'h2632] <= 8'h29;
		memory[16'h2633] <= 8'h1a;
		memory[16'h2634] <= 8'hc0;
		memory[16'h2635] <= 8'h3a;
		memory[16'h2636] <= 8'h40;
		memory[16'h2637] <= 8'h18;
		memory[16'h2638] <= 8'h5;
		memory[16'h2639] <= 8'h50;
		memory[16'h263a] <= 8'he0;
		memory[16'h263b] <= 8'h4f;
		memory[16'h263c] <= 8'h78;
		memory[16'h263d] <= 8'hf2;
		memory[16'h263e] <= 8'h3d;
		memory[16'h263f] <= 8'h3f;
		memory[16'h2640] <= 8'hf0;
		memory[16'h2641] <= 8'h1b;
		memory[16'h2642] <= 8'h66;
		memory[16'h2643] <= 8'h97;
		memory[16'h2644] <= 8'h6a;
		memory[16'h2645] <= 8'hb1;
		memory[16'h2646] <= 8'he;
		memory[16'h2647] <= 8'h84;
		memory[16'h2648] <= 8'h84;
		memory[16'h2649] <= 8'he2;
		memory[16'h264a] <= 8'h62;
		memory[16'h264b] <= 8'hfa;
		memory[16'h264c] <= 8'h37;
		memory[16'h264d] <= 8'h23;
		memory[16'h264e] <= 8'ha7;
		memory[16'h264f] <= 8'h94;
		memory[16'h2650] <= 8'hb5;
		memory[16'h2651] <= 8'hd0;
		memory[16'h2652] <= 8'hae;
		memory[16'h2653] <= 8'h75;
		memory[16'h2654] <= 8'ha;
		memory[16'h2655] <= 8'hee;
		memory[16'h2656] <= 8'h8d;
		memory[16'h2657] <= 8'hf;
		memory[16'h2658] <= 8'h3e;
		memory[16'h2659] <= 8'h6d;
		memory[16'h265a] <= 8'h5f;
		memory[16'h265b] <= 8'hb6;
		memory[16'h265c] <= 8'h60;
		memory[16'h265d] <= 8'h9c;
		memory[16'h265e] <= 8'hf5;
		memory[16'h265f] <= 8'h50;
		memory[16'h2660] <= 8'hb7;
		memory[16'h2661] <= 8'h5c;
		memory[16'h2662] <= 8'he7;
		memory[16'h2663] <= 8'h21;
		memory[16'h2664] <= 8'hd;
		memory[16'h2665] <= 8'hf6;
		memory[16'h2666] <= 8'ha5;
		memory[16'h2667] <= 8'h91;
		memory[16'h2668] <= 8'hd8;
		memory[16'h2669] <= 8'h8;
		memory[16'h266a] <= 8'h8b;
		memory[16'h266b] <= 8'h10;
		memory[16'h266c] <= 8'h2b;
		memory[16'h266d] <= 8'h32;
		memory[16'h266e] <= 8'ha4;
		memory[16'h266f] <= 8'he0;
		memory[16'h2670] <= 8'h2;
		memory[16'h2671] <= 8'h52;
		memory[16'h2672] <= 8'h55;
		memory[16'h2673] <= 8'hc;
		memory[16'h2674] <= 8'h40;
		memory[16'h2675] <= 8'he2;
		memory[16'h2676] <= 8'h1c;
		memory[16'h2677] <= 8'h7f;
		memory[16'h2678] <= 8'h50;
		memory[16'h2679] <= 8'h7b;
		memory[16'h267a] <= 8'h35;
		memory[16'h267b] <= 8'hb0;
		memory[16'h267c] <= 8'h17;
		memory[16'h267d] <= 8'h2b;
		memory[16'h267e] <= 8'h0;
		memory[16'h267f] <= 8'hce;
		memory[16'h2680] <= 8'h87;
		memory[16'h2681] <= 8'he8;
		memory[16'h2682] <= 8'hef;
		memory[16'h2683] <= 8'h94;
		memory[16'h2684] <= 8'hde;
		memory[16'h2685] <= 8'h94;
		memory[16'h2686] <= 8'h25;
		memory[16'h2687] <= 8'hb6;
		memory[16'h2688] <= 8'h9c;
		memory[16'h2689] <= 8'hb0;
		memory[16'h268a] <= 8'hc6;
		memory[16'h268b] <= 8'hc8;
		memory[16'h268c] <= 8'he3;
		memory[16'h268d] <= 8'h6a;
		memory[16'h268e] <= 8'ha8;
		memory[16'h268f] <= 8'he5;
		memory[16'h2690] <= 8'hbc;
		memory[16'h2691] <= 8'hfe;
		memory[16'h2692] <= 8'hf2;
		memory[16'h2693] <= 8'hfd;
		memory[16'h2694] <= 8'he0;
		memory[16'h2695] <= 8'he;
		memory[16'h2696] <= 8'h7c;
		memory[16'h2697] <= 8'h30;
		memory[16'h2698] <= 8'h89;
		memory[16'h2699] <= 8'hb1;
		memory[16'h269a] <= 8'he0;
		memory[16'h269b] <= 8'ha0;
		memory[16'h269c] <= 8'hdc;
		memory[16'h269d] <= 8'he1;
		memory[16'h269e] <= 8'h6e;
		memory[16'h269f] <= 8'h63;
		memory[16'h26a0] <= 8'hc9;
		memory[16'h26a1] <= 8'h5d;
		memory[16'h26a2] <= 8'hf7;
		memory[16'h26a3] <= 8'ha7;
		memory[16'h26a4] <= 8'hf1;
		memory[16'h26a5] <= 8'h1c;
		memory[16'h26a6] <= 8'h5d;
		memory[16'h26a7] <= 8'h8e;
		memory[16'h26a8] <= 8'hcd;
		memory[16'h26a9] <= 8'h24;
		memory[16'h26aa] <= 8'h56;
		memory[16'h26ab] <= 8'hb0;
		memory[16'h26ac] <= 8'h8e;
		memory[16'h26ad] <= 8'hfe;
		memory[16'h26ae] <= 8'h95;
		memory[16'h26af] <= 8'h4b;
		memory[16'h26b0] <= 8'hfc;
		memory[16'h26b1] <= 8'h87;
		memory[16'h26b2] <= 8'h48;
		memory[16'h26b3] <= 8'hdd;
		memory[16'h26b4] <= 8'h95;
		memory[16'h26b5] <= 8'hc4;
		memory[16'h26b6] <= 8'hd;
		memory[16'h26b7] <= 8'h1e;
		memory[16'h26b8] <= 8'h75;
		memory[16'h26b9] <= 8'hee;
		memory[16'h26ba] <= 8'hbe;
		memory[16'h26bb] <= 8'h52;
		memory[16'h26bc] <= 8'hcf;
		memory[16'h26bd] <= 8'h2c;
		memory[16'h26be] <= 8'hb5;
		memory[16'h26bf] <= 8'h98;
		memory[16'h26c0] <= 8'h89;
		memory[16'h26c1] <= 8'had;
		memory[16'h26c2] <= 8'h3f;
		memory[16'h26c3] <= 8'h7b;
		memory[16'h26c4] <= 8'hc9;
		memory[16'h26c5] <= 8'h9c;
		memory[16'h26c6] <= 8'h9;
		memory[16'h26c7] <= 8'h96;
		memory[16'h26c8] <= 8'hc0;
		memory[16'h26c9] <= 8'h5f;
		memory[16'h26ca] <= 8'h46;
		memory[16'h26cb] <= 8'h4f;
		memory[16'h26cc] <= 8'h5d;
		memory[16'h26cd] <= 8'hdc;
		memory[16'h26ce] <= 8'h9a;
		memory[16'h26cf] <= 8'h5a;
		memory[16'h26d0] <= 8'h63;
		memory[16'h26d1] <= 8'he2;
		memory[16'h26d2] <= 8'h37;
		memory[16'h26d3] <= 8'hf9;
		memory[16'h26d4] <= 8'ha6;
		memory[16'h26d5] <= 8'h44;
		memory[16'h26d6] <= 8'h17;
		memory[16'h26d7] <= 8'h1b;
		memory[16'h26d8] <= 8'h32;
		memory[16'h26d9] <= 8'hd6;
		memory[16'h26da] <= 8'h6d;
		memory[16'h26db] <= 8'h1;
		memory[16'h26dc] <= 8'h2;
		memory[16'h26dd] <= 8'h23;
		memory[16'h26de] <= 8'h99;
		memory[16'h26df] <= 8'h8c;
		memory[16'h26e0] <= 8'hd0;
		memory[16'h26e1] <= 8'hd8;
		memory[16'h26e2] <= 8'h7;
		memory[16'h26e3] <= 8'h99;
		memory[16'h26e4] <= 8'h75;
		memory[16'h26e5] <= 8'h10;
		memory[16'h26e6] <= 8'h30;
		memory[16'h26e7] <= 8'h35;
		memory[16'h26e8] <= 8'h6f;
		memory[16'h26e9] <= 8'h76;
		memory[16'h26ea] <= 8'h84;
		memory[16'h26eb] <= 8'hcc;
		memory[16'h26ec] <= 8'h52;
		memory[16'h26ed] <= 8'h1e;
		memory[16'h26ee] <= 8'h26;
		memory[16'h26ef] <= 8'hb6;
		memory[16'h26f0] <= 8'h0;
		memory[16'h26f1] <= 8'h5d;
		memory[16'h26f2] <= 8'haf;
		memory[16'h26f3] <= 8'ha6;
		memory[16'h26f4] <= 8'ha2;
		memory[16'h26f5] <= 8'hc6;
		memory[16'h26f6] <= 8'hc2;
		memory[16'h26f7] <= 8'hd4;
		memory[16'h26f8] <= 8'h9c;
		memory[16'h26f9] <= 8'h2f;
		memory[16'h26fa] <= 8'hd6;
		memory[16'h26fb] <= 8'h9f;
		memory[16'h26fc] <= 8'h52;
		memory[16'h26fd] <= 8'h6f;
		memory[16'h26fe] <= 8'h2b;
		memory[16'h26ff] <= 8'h22;
		memory[16'h2700] <= 8'h48;
		memory[16'h2701] <= 8'h32;
		memory[16'h2702] <= 8'hbc;
		memory[16'h2703] <= 8'hbd;
		memory[16'h2704] <= 8'h42;
		memory[16'h2705] <= 8'hec;
		memory[16'h2706] <= 8'hf2;
		memory[16'h2707] <= 8'hb1;
		memory[16'h2708] <= 8'h62;
		memory[16'h2709] <= 8'h77;
		memory[16'h270a] <= 8'h7d;
		memory[16'h270b] <= 8'hb5;
		memory[16'h270c] <= 8'h95;
		memory[16'h270d] <= 8'ha4;
		memory[16'h270e] <= 8'h6b;
		memory[16'h270f] <= 8'h96;
		memory[16'h2710] <= 8'h1;
		memory[16'h2711] <= 8'h1a;
		memory[16'h2712] <= 8'h3c;
		memory[16'h2713] <= 8'ha3;
		memory[16'h2714] <= 8'he0;
		memory[16'h2715] <= 8'hfe;
		memory[16'h2716] <= 8'h78;
		memory[16'h2717] <= 8'h7d;
		memory[16'h2718] <= 8'h2e;
		memory[16'h2719] <= 8'h4e;
		memory[16'h271a] <= 8'h1c;
		memory[16'h271b] <= 8'h80;
		memory[16'h271c] <= 8'hbd;
		memory[16'h271d] <= 8'h47;
		memory[16'h271e] <= 8'ha3;
		memory[16'h271f] <= 8'h5;
		memory[16'h2720] <= 8'h79;
		memory[16'h2721] <= 8'h5f;
		memory[16'h2722] <= 8'hc2;
		memory[16'h2723] <= 8'hbb;
		memory[16'h2724] <= 8'h4b;
		memory[16'h2725] <= 8'hb5;
		memory[16'h2726] <= 8'h6c;
		memory[16'h2727] <= 8'had;
		memory[16'h2728] <= 8'h2c;
		memory[16'h2729] <= 8'he9;
		memory[16'h272a] <= 8'h62;
		memory[16'h272b] <= 8'hc1;
		memory[16'h272c] <= 8'h8d;
		memory[16'h272d] <= 8'hcd;
		memory[16'h272e] <= 8'h57;
		memory[16'h272f] <= 8'h8f;
		memory[16'h2730] <= 8'he7;
		memory[16'h2731] <= 8'h94;
		memory[16'h2732] <= 8'h32;
		memory[16'h2733] <= 8'hc8;
		memory[16'h2734] <= 8'h92;
		memory[16'h2735] <= 8'haa;
		memory[16'h2736] <= 8'h45;
		memory[16'h2737] <= 8'hc0;
		memory[16'h2738] <= 8'hf8;
		memory[16'h2739] <= 8'h61;
		memory[16'h273a] <= 8'h41;
		memory[16'h273b] <= 8'hb6;
		memory[16'h273c] <= 8'ha8;
		memory[16'h273d] <= 8'he4;
		memory[16'h273e] <= 8'hbb;
		memory[16'h273f] <= 8'h21;
		memory[16'h2740] <= 8'h43;
		memory[16'h2741] <= 8'h7e;
		memory[16'h2742] <= 8'hdc;
		memory[16'h2743] <= 8'h8e;
		memory[16'h2744] <= 8'h33;
		memory[16'h2745] <= 8'h48;
		memory[16'h2746] <= 8'h3b;
		memory[16'h2747] <= 8'h5f;
		memory[16'h2748] <= 8'h31;
		memory[16'h2749] <= 8'h9e;
		memory[16'h274a] <= 8'h20;
		memory[16'h274b] <= 8'hbf;
		memory[16'h274c] <= 8'h6b;
		memory[16'h274d] <= 8'h78;
		memory[16'h274e] <= 8'h4e;
		memory[16'h274f] <= 8'h53;
		memory[16'h2750] <= 8'hc;
		memory[16'h2751] <= 8'h80;
		memory[16'h2752] <= 8'h1b;
		memory[16'h2753] <= 8'h9e;
		memory[16'h2754] <= 8'h2b;
		memory[16'h2755] <= 8'h60;
		memory[16'h2756] <= 8'h5f;
		memory[16'h2757] <= 8'h23;
		memory[16'h2758] <= 8'hc1;
		memory[16'h2759] <= 8'ha0;
		memory[16'h275a] <= 8'hd9;
		memory[16'h275b] <= 8'h69;
		memory[16'h275c] <= 8'h84;
		memory[16'h275d] <= 8'h95;
		memory[16'h275e] <= 8'h8a;
		memory[16'h275f] <= 8'hc7;
		memory[16'h2760] <= 8'h13;
		memory[16'h2761] <= 8'h66;
		memory[16'h2762] <= 8'h55;
		memory[16'h2763] <= 8'h46;
		memory[16'h2764] <= 8'hae;
		memory[16'h2765] <= 8'h90;
		memory[16'h2766] <= 8'ha5;
		memory[16'h2767] <= 8'hdf;
		memory[16'h2768] <= 8'h2e;
		memory[16'h2769] <= 8'hc5;
		memory[16'h276a] <= 8'h9e;
		memory[16'h276b] <= 8'h9a;
		memory[16'h276c] <= 8'h3d;
		memory[16'h276d] <= 8'hec;
		memory[16'h276e] <= 8'hed;
		memory[16'h276f] <= 8'h49;
		memory[16'h2770] <= 8'h6d;
		memory[16'h2771] <= 8'h8;
		memory[16'h2772] <= 8'he8;
		memory[16'h2773] <= 8'h98;
		memory[16'h2774] <= 8'h68;
		memory[16'h2775] <= 8'h47;
		memory[16'h2776] <= 8'hbb;
		memory[16'h2777] <= 8'h29;
		memory[16'h2778] <= 8'he7;
		memory[16'h2779] <= 8'h95;
		memory[16'h277a] <= 8'h92;
		memory[16'h277b] <= 8'h6b;
		memory[16'h277c] <= 8'h2a;
		memory[16'h277d] <= 8'h1c;
		memory[16'h277e] <= 8'h32;
		memory[16'h277f] <= 8'h3d;
		memory[16'h2780] <= 8'h82;
		memory[16'h2781] <= 8'h87;
		memory[16'h2782] <= 8'h83;
		memory[16'h2783] <= 8'h30;
		memory[16'h2784] <= 8'h17;
		memory[16'h2785] <= 8'h28;
		memory[16'h2786] <= 8'hf;
		memory[16'h2787] <= 8'h46;
		memory[16'h2788] <= 8'hed;
		memory[16'h2789] <= 8'hae;
		memory[16'h278a] <= 8'he0;
		memory[16'h278b] <= 8'h2b;
		memory[16'h278c] <= 8'h9a;
		memory[16'h278d] <= 8'hcd;
		memory[16'h278e] <= 8'h74;
		memory[16'h278f] <= 8'h7;
		memory[16'h2790] <= 8'hd5;
		memory[16'h2791] <= 8'h5c;
		memory[16'h2792] <= 8'h9f;
		memory[16'h2793] <= 8'h3d;
		memory[16'h2794] <= 8'ha3;
		memory[16'h2795] <= 8'h5b;
		memory[16'h2796] <= 8'h66;
		memory[16'h2797] <= 8'h8a;
		memory[16'h2798] <= 8'hf0;
		memory[16'h2799] <= 8'hf8;
		memory[16'h279a] <= 8'hf5;
		memory[16'h279b] <= 8'h1a;
		memory[16'h279c] <= 8'h14;
		memory[16'h279d] <= 8'h27;
		memory[16'h279e] <= 8'h57;
		memory[16'h279f] <= 8'h96;
		memory[16'h27a0] <= 8'hae;
		memory[16'h27a1] <= 8'hda;
		memory[16'h27a2] <= 8'hc6;
		memory[16'h27a3] <= 8'hc6;
		memory[16'h27a4] <= 8'h2;
		memory[16'h27a5] <= 8'hd5;
		memory[16'h27a6] <= 8'hc;
		memory[16'h27a7] <= 8'hef;
		memory[16'h27a8] <= 8'h83;
		memory[16'h27a9] <= 8'hec;
		memory[16'h27aa] <= 8'h1a;
		memory[16'h27ab] <= 8'h1e;
		memory[16'h27ac] <= 8'hb9;
		memory[16'h27ad] <= 8'h8f;
		memory[16'h27ae] <= 8'h25;
		memory[16'h27af] <= 8'h8e;
		memory[16'h27b0] <= 8'heb;
		memory[16'h27b1] <= 8'hc5;
		memory[16'h27b2] <= 8'hcb;
		memory[16'h27b3] <= 8'h8f;
		memory[16'h27b4] <= 8'h20;
		memory[16'h27b5] <= 8'h31;
		memory[16'h27b6] <= 8'h19;
		memory[16'h27b7] <= 8'h10;
		memory[16'h27b8] <= 8'h29;
		memory[16'h27b9] <= 8'hf;
		memory[16'h27ba] <= 8'h2a;
		memory[16'h27bb] <= 8'h3d;
		memory[16'h27bc] <= 8'h36;
		memory[16'h27bd] <= 8'h81;
		memory[16'h27be] <= 8'hd3;
		memory[16'h27bf] <= 8'he5;
		memory[16'h27c0] <= 8'h5b;
		memory[16'h27c1] <= 8'h99;
		memory[16'h27c2] <= 8'hab;
		memory[16'h27c3] <= 8'h5d;
		memory[16'h27c4] <= 8'h6e;
		memory[16'h27c5] <= 8'hb7;
		memory[16'h27c6] <= 8'h4c;
		memory[16'h27c7] <= 8'hf2;
		memory[16'h27c8] <= 8'ha3;
		memory[16'h27c9] <= 8'h67;
		memory[16'h27ca] <= 8'h10;
		memory[16'h27cb] <= 8'h5c;
		memory[16'h27cc] <= 8'hf6;
		memory[16'h27cd] <= 8'h35;
		memory[16'h27ce] <= 8'hea;
		memory[16'h27cf] <= 8'he1;
		memory[16'h27d0] <= 8'hfa;
		memory[16'h27d1] <= 8'hb5;
		memory[16'h27d2] <= 8'h70;
		memory[16'h27d3] <= 8'h1a;
		memory[16'h27d4] <= 8'he6;
		memory[16'h27d5] <= 8'h8a;
		memory[16'h27d6] <= 8'h2a;
		memory[16'h27d7] <= 8'hf;
		memory[16'h27d8] <= 8'h99;
		memory[16'h27d9] <= 8'h54;
		memory[16'h27da] <= 8'h4c;
		memory[16'h27db] <= 8'hcf;
		memory[16'h27dc] <= 8'hd5;
		memory[16'h27dd] <= 8'h1f;
		memory[16'h27de] <= 8'hb4;
		memory[16'h27df] <= 8'h30;
		memory[16'h27e0] <= 8'hb8;
		memory[16'h27e1] <= 8'h5f;
		memory[16'h27e2] <= 8'h8d;
		memory[16'h27e3] <= 8'h26;
		memory[16'h27e4] <= 8'h16;
		memory[16'h27e5] <= 8'hda;
		memory[16'h27e6] <= 8'h18;
		memory[16'h27e7] <= 8'hb9;
		memory[16'h27e8] <= 8'h41;
		memory[16'h27e9] <= 8'h28;
		memory[16'h27ea] <= 8'h15;
		memory[16'h27eb] <= 8'h37;
		memory[16'h27ec] <= 8'h5e;
		memory[16'h27ed] <= 8'hff;
		memory[16'h27ee] <= 8'h18;
		memory[16'h27ef] <= 8'h58;
		memory[16'h27f0] <= 8'hb4;
		memory[16'h27f1] <= 8'h89;
		memory[16'h27f2] <= 8'h73;
		memory[16'h27f3] <= 8'h9a;
		memory[16'h27f4] <= 8'h13;
		memory[16'h27f5] <= 8'h9d;
		memory[16'h27f6] <= 8'ha9;
		memory[16'h27f7] <= 8'hac;
		memory[16'h27f8] <= 8'hf2;
		memory[16'h27f9] <= 8'hf5;
		memory[16'h27fa] <= 8'h7b;
		memory[16'h27fb] <= 8'hc7;
		memory[16'h27fc] <= 8'h14;
		memory[16'h27fd] <= 8'h30;
		memory[16'h27fe] <= 8'hf8;
		memory[16'h27ff] <= 8'hcc;
		memory[16'h2800] <= 8'h8f;
		memory[16'h2801] <= 8'h85;
		memory[16'h2802] <= 8'hf3;
		memory[16'h2803] <= 8'ha6;
		memory[16'h2804] <= 8'h5f;
		memory[16'h2805] <= 8'hb;
		memory[16'h2806] <= 8'h5f;
		memory[16'h2807] <= 8'ha0;
		memory[16'h2808] <= 8'h34;
		memory[16'h2809] <= 8'h75;
		memory[16'h280a] <= 8'hd7;
		memory[16'h280b] <= 8'h92;
		memory[16'h280c] <= 8'h74;
		memory[16'h280d] <= 8'hf0;
		memory[16'h280e] <= 8'hea;
		memory[16'h280f] <= 8'h29;
		memory[16'h2810] <= 8'h79;
		memory[16'h2811] <= 8'h5d;
		memory[16'h2812] <= 8'hc3;
		memory[16'h2813] <= 8'h8c;
		memory[16'h2814] <= 8'hfb;
		memory[16'h2815] <= 8'h6d;
		memory[16'h2816] <= 8'h38;
		memory[16'h2817] <= 8'hed;
		memory[16'h2818] <= 8'h62;
		memory[16'h2819] <= 8'hb3;
		memory[16'h281a] <= 8'hb4;
		memory[16'h281b] <= 8'h77;
		memory[16'h281c] <= 8'he3;
		memory[16'h281d] <= 8'hac;
		memory[16'h281e] <= 8'h43;
		memory[16'h281f] <= 8'h73;
		memory[16'h2820] <= 8'h32;
		memory[16'h2821] <= 8'h36;
		memory[16'h2822] <= 8'h19;
		memory[16'h2823] <= 8'h91;
		memory[16'h2824] <= 8'h42;
		memory[16'h2825] <= 8'h78;
		memory[16'h2826] <= 8'h32;
		memory[16'h2827] <= 8'h76;
		memory[16'h2828] <= 8'hed;
		memory[16'h2829] <= 8'h9;
		memory[16'h282a] <= 8'h8;
		memory[16'h282b] <= 8'h62;
		memory[16'h282c] <= 8'hf9;
		memory[16'h282d] <= 8'hf2;
		memory[16'h282e] <= 8'h8b;
		memory[16'h282f] <= 8'h72;
		memory[16'h2830] <= 8'h50;
		memory[16'h2831] <= 8'h4e;
		memory[16'h2832] <= 8'hfe;
		memory[16'h2833] <= 8'h4b;
		memory[16'h2834] <= 8'hbb;
		memory[16'h2835] <= 8'h36;
		memory[16'h2836] <= 8'h38;
		memory[16'h2837] <= 8'h1e;
		memory[16'h2838] <= 8'hea;
		memory[16'h2839] <= 8'hec;
		memory[16'h283a] <= 8'h95;
		memory[16'h283b] <= 8'hcd;
		memory[16'h283c] <= 8'h99;
		memory[16'h283d] <= 8'hd8;
		memory[16'h283e] <= 8'h40;
		memory[16'h283f] <= 8'hcb;
		memory[16'h2840] <= 8'hf;
		memory[16'h2841] <= 8'h59;
		memory[16'h2842] <= 8'h5c;
		memory[16'h2843] <= 8'h51;
		memory[16'h2844] <= 8'hd2;
		memory[16'h2845] <= 8'h8e;
		memory[16'h2846] <= 8'hc7;
		memory[16'h2847] <= 8'hbf;
		memory[16'h2848] <= 8'h98;
		memory[16'h2849] <= 8'hcf;
		memory[16'h284a] <= 8'h21;
		memory[16'h284b] <= 8'h91;
		memory[16'h284c] <= 8'hc1;
		memory[16'h284d] <= 8'hac;
		memory[16'h284e] <= 8'h4;
		memory[16'h284f] <= 8'h11;
		memory[16'h2850] <= 8'hfb;
		memory[16'h2851] <= 8'h2;
		memory[16'h2852] <= 8'h5c;
		memory[16'h2853] <= 8'hb6;
		memory[16'h2854] <= 8'h39;
		memory[16'h2855] <= 8'h94;
		memory[16'h2856] <= 8'hd4;
		memory[16'h2857] <= 8'h23;
		memory[16'h2858] <= 8'h81;
		memory[16'h2859] <= 8'h69;
		memory[16'h285a] <= 8'hf0;
		memory[16'h285b] <= 8'h1a;
		memory[16'h285c] <= 8'h42;
		memory[16'h285d] <= 8'h31;
		memory[16'h285e] <= 8'he5;
		memory[16'h285f] <= 8'h51;
		memory[16'h2860] <= 8'h8a;
		memory[16'h2861] <= 8'h41;
		memory[16'h2862] <= 8'ha2;
		memory[16'h2863] <= 8'h5c;
		memory[16'h2864] <= 8'hd0;
		memory[16'h2865] <= 8'h69;
		memory[16'h2866] <= 8'h1c;
		memory[16'h2867] <= 8'h68;
		memory[16'h2868] <= 8'h38;
		memory[16'h2869] <= 8'h3d;
		memory[16'h286a] <= 8'hf9;
		memory[16'h286b] <= 8'hf9;
		memory[16'h286c] <= 8'hea;
		memory[16'h286d] <= 8'hfd;
		memory[16'h286e] <= 8'hb;
		memory[16'h286f] <= 8'he5;
		memory[16'h2870] <= 8'h0;
		memory[16'h2871] <= 8'h67;
		memory[16'h2872] <= 8'h9b;
		memory[16'h2873] <= 8'h39;
		memory[16'h2874] <= 8'hfc;
		memory[16'h2875] <= 8'h70;
		memory[16'h2876] <= 8'h5c;
		memory[16'h2877] <= 8'h7d;
		memory[16'h2878] <= 8'hd9;
		memory[16'h2879] <= 8'h4c;
		memory[16'h287a] <= 8'h97;
		memory[16'h287b] <= 8'h1b;
		memory[16'h287c] <= 8'h7d;
		memory[16'h287d] <= 8'h7c;
		memory[16'h287e] <= 8'h6c;
		memory[16'h287f] <= 8'h8;
		memory[16'h2880] <= 8'hbd;
		memory[16'h2881] <= 8'he;
		memory[16'h2882] <= 8'h64;
		memory[16'h2883] <= 8'h8d;
		memory[16'h2884] <= 8'h77;
		memory[16'h2885] <= 8'h80;
		memory[16'h2886] <= 8'hf5;
		memory[16'h2887] <= 8'haf;
		memory[16'h2888] <= 8'hbe;
		memory[16'h2889] <= 8'hef;
		memory[16'h288a] <= 8'ha9;
		memory[16'h288b] <= 8'ha8;
		memory[16'h288c] <= 8'hec;
		memory[16'h288d] <= 8'hb4;
		memory[16'h288e] <= 8'h8d;
		memory[16'h288f] <= 8'hec;
		memory[16'h2890] <= 8'h1b;
		memory[16'h2891] <= 8'h28;
		memory[16'h2892] <= 8'h25;
		memory[16'h2893] <= 8'h17;
		memory[16'h2894] <= 8'h98;
		memory[16'h2895] <= 8'h81;
		memory[16'h2896] <= 8'h94;
		memory[16'h2897] <= 8'h72;
		memory[16'h2898] <= 8'hce;
		memory[16'h2899] <= 8'h2b;
		memory[16'h289a] <= 8'h8d;
		memory[16'h289b] <= 8'h4b;
		memory[16'h289c] <= 8'ha7;
		memory[16'h289d] <= 8'hfa;
		memory[16'h289e] <= 8'h53;
		memory[16'h289f] <= 8'h65;
		memory[16'h28a0] <= 8'h8;
		memory[16'h28a1] <= 8'hb8;
		memory[16'h28a2] <= 8'hf2;
		memory[16'h28a3] <= 8'h80;
		memory[16'h28a4] <= 8'h38;
		memory[16'h28a5] <= 8'he8;
		memory[16'h28a6] <= 8'h2f;
		memory[16'h28a7] <= 8'hf6;
		memory[16'h28a8] <= 8'hd7;
		memory[16'h28a9] <= 8'hd8;
		memory[16'h28aa] <= 8'h9e;
		memory[16'h28ab] <= 8'hc3;
		memory[16'h28ac] <= 8'h8c;
		memory[16'h28ad] <= 8'h2b;
		memory[16'h28ae] <= 8'hb0;
		memory[16'h28af] <= 8'ha8;
		memory[16'h28b0] <= 8'h54;
		memory[16'h28b1] <= 8'hd5;
		memory[16'h28b2] <= 8'hbf;
		memory[16'h28b3] <= 8'hec;
		memory[16'h28b4] <= 8'h57;
		memory[16'h28b5] <= 8'h54;
		memory[16'h28b6] <= 8'h5e;
		memory[16'h28b7] <= 8'h25;
		memory[16'h28b8] <= 8'h7f;
		memory[16'h28b9] <= 8'hec;
		memory[16'h28ba] <= 8'h70;
		memory[16'h28bb] <= 8'h27;
		memory[16'h28bc] <= 8'he6;
		memory[16'h28bd] <= 8'hc4;
		memory[16'h28be] <= 8'h8c;
		memory[16'h28bf] <= 8'hee;
		memory[16'h28c0] <= 8'h7c;
		memory[16'h28c1] <= 8'h7e;
		memory[16'h28c2] <= 8'h6e;
		memory[16'h28c3] <= 8'hb4;
		memory[16'h28c4] <= 8'h66;
		memory[16'h28c5] <= 8'h9e;
		memory[16'h28c6] <= 8'hab;
		memory[16'h28c7] <= 8'h3d;
		memory[16'h28c8] <= 8'h76;
		memory[16'h28c9] <= 8'h49;
		memory[16'h28ca] <= 8'h1;
		memory[16'h28cb] <= 8'h3;
		memory[16'h28cc] <= 8'h75;
		memory[16'h28cd] <= 8'hb1;
		memory[16'h28ce] <= 8'hab;
		memory[16'h28cf] <= 8'hc9;
		memory[16'h28d0] <= 8'h86;
		memory[16'h28d1] <= 8'h6a;
		memory[16'h28d2] <= 8'hb5;
		memory[16'h28d3] <= 8'hdd;
		memory[16'h28d4] <= 8'hbe;
		memory[16'h28d5] <= 8'h14;
		memory[16'h28d6] <= 8'h2;
		memory[16'h28d7] <= 8'h3e;
		memory[16'h28d8] <= 8'h0;
		memory[16'h28d9] <= 8'h73;
		memory[16'h28da] <= 8'h65;
		memory[16'h28db] <= 8'he6;
		memory[16'h28dc] <= 8'h37;
		memory[16'h28dd] <= 8'hf1;
		memory[16'h28de] <= 8'hd4;
		memory[16'h28df] <= 8'hb3;
		memory[16'h28e0] <= 8'h6f;
		memory[16'h28e1] <= 8'h43;
		memory[16'h28e2] <= 8'h67;
		memory[16'h28e3] <= 8'hd6;
		memory[16'h28e4] <= 8'he1;
		memory[16'h28e5] <= 8'h12;
		memory[16'h28e6] <= 8'h13;
		memory[16'h28e7] <= 8'h57;
		memory[16'h28e8] <= 8'h5c;
		memory[16'h28e9] <= 8'h14;
		memory[16'h28ea] <= 8'h5a;
		memory[16'h28eb] <= 8'hd1;
		memory[16'h28ec] <= 8'hc5;
		memory[16'h28ed] <= 8'h5;
		memory[16'h28ee] <= 8'h9a;
		memory[16'h28ef] <= 8'h4c;
		memory[16'h28f0] <= 8'h70;
		memory[16'h28f1] <= 8'h4f;
		memory[16'h28f2] <= 8'h29;
		memory[16'h28f3] <= 8'h2e;
		memory[16'h28f4] <= 8'h63;
		memory[16'h28f5] <= 8'h2c;
		memory[16'h28f6] <= 8'h6c;
		memory[16'h28f7] <= 8'h63;
		memory[16'h28f8] <= 8'h9f;
		memory[16'h28f9] <= 8'hd1;
		memory[16'h28fa] <= 8'h49;
		memory[16'h28fb] <= 8'hd6;
		memory[16'h28fc] <= 8'hc2;
		memory[16'h28fd] <= 8'h1e;
		memory[16'h28fe] <= 8'h89;
		memory[16'h28ff] <= 8'h32;
		memory[16'h2900] <= 8'h61;
		memory[16'h2901] <= 8'hf0;
		memory[16'h2902] <= 8'h8;
		memory[16'h2903] <= 8'h42;
		memory[16'h2904] <= 8'h3;
		memory[16'h2905] <= 8'h1b;
		memory[16'h2906] <= 8'h99;
		memory[16'h2907] <= 8'h5f;
		memory[16'h2908] <= 8'h30;
		memory[16'h2909] <= 8'hf4;
		memory[16'h290a] <= 8'h30;
		memory[16'h290b] <= 8'hf5;
		memory[16'h290c] <= 8'hf9;
		memory[16'h290d] <= 8'hca;
		memory[16'h290e] <= 8'h41;
		memory[16'h290f] <= 8'h69;
		memory[16'h2910] <= 8'h19;
		memory[16'h2911] <= 8'h6b;
		memory[16'h2912] <= 8'h98;
		memory[16'h2913] <= 8'h7d;
		memory[16'h2914] <= 8'h97;
		memory[16'h2915] <= 8'h4;
		memory[16'h2916] <= 8'he0;
		memory[16'h2917] <= 8'h36;
		memory[16'h2918] <= 8'hd6;
		memory[16'h2919] <= 8'h2a;
		memory[16'h291a] <= 8'hc;
		memory[16'h291b] <= 8'h98;
		memory[16'h291c] <= 8'h48;
		memory[16'h291d] <= 8'h95;
		memory[16'h291e] <= 8'hca;
		memory[16'h291f] <= 8'ha9;
		memory[16'h2920] <= 8'h85;
		memory[16'h2921] <= 8'hd2;
		memory[16'h2922] <= 8'heb;
		memory[16'h2923] <= 8'h88;
		memory[16'h2924] <= 8'hee;
		memory[16'h2925] <= 8'h84;
		memory[16'h2926] <= 8'he7;
		memory[16'h2927] <= 8'h1e;
		memory[16'h2928] <= 8'h78;
		memory[16'h2929] <= 8'h17;
		memory[16'h292a] <= 8'h13;
		memory[16'h292b] <= 8'h72;
		memory[16'h292c] <= 8'he1;
		memory[16'h292d] <= 8'h55;
		memory[16'h292e] <= 8'hdb;
		memory[16'h292f] <= 8'hfb;
		memory[16'h2930] <= 8'hc0;
		memory[16'h2931] <= 8'h73;
		memory[16'h2932] <= 8'h78;
		memory[16'h2933] <= 8'h57;
		memory[16'h2934] <= 8'h78;
		memory[16'h2935] <= 8'h58;
		memory[16'h2936] <= 8'h8d;
		memory[16'h2937] <= 8'h4e;
		memory[16'h2938] <= 8'h82;
		memory[16'h2939] <= 8'h99;
		memory[16'h293a] <= 8'he6;
		memory[16'h293b] <= 8'hca;
		memory[16'h293c] <= 8'h2e;
		memory[16'h293d] <= 8'hb1;
		memory[16'h293e] <= 8'h73;
		memory[16'h293f] <= 8'hb3;
		memory[16'h2940] <= 8'h83;
		memory[16'h2941] <= 8'h5e;
		memory[16'h2942] <= 8'h3c;
		memory[16'h2943] <= 8'h71;
		memory[16'h2944] <= 8'he3;
		memory[16'h2945] <= 8'h23;
		memory[16'h2946] <= 8'h8f;
		memory[16'h2947] <= 8'h5b;
		memory[16'h2948] <= 8'h3b;
		memory[16'h2949] <= 8'ha3;
		memory[16'h294a] <= 8'hcd;
		memory[16'h294b] <= 8'h1c;
		memory[16'h294c] <= 8'hf8;
		memory[16'h294d] <= 8'ha9;
		memory[16'h294e] <= 8'h17;
		memory[16'h294f] <= 8'hb8;
		memory[16'h2950] <= 8'h1c;
		memory[16'h2951] <= 8'h8f;
		memory[16'h2952] <= 8'hf;
		memory[16'h2953] <= 8'h94;
		memory[16'h2954] <= 8'he8;
		memory[16'h2955] <= 8'h9c;
		memory[16'h2956] <= 8'he2;
		memory[16'h2957] <= 8'h6a;
		memory[16'h2958] <= 8'h35;
		memory[16'h2959] <= 8'hc9;
		memory[16'h295a] <= 8'h35;
		memory[16'h295b] <= 8'h63;
		memory[16'h295c] <= 8'h7a;
		memory[16'h295d] <= 8'ha8;
		memory[16'h295e] <= 8'h16;
		memory[16'h295f] <= 8'hfd;
		memory[16'h2960] <= 8'h7;
		memory[16'h2961] <= 8'h52;
		memory[16'h2962] <= 8'h6f;
		memory[16'h2963] <= 8'hea;
		memory[16'h2964] <= 8'h76;
		memory[16'h2965] <= 8'hfe;
		memory[16'h2966] <= 8'h45;
		memory[16'h2967] <= 8'hb1;
		memory[16'h2968] <= 8'ha1;
		memory[16'h2969] <= 8'h13;
		memory[16'h296a] <= 8'hcd;
		memory[16'h296b] <= 8'h99;
		memory[16'h296c] <= 8'hbc;
		memory[16'h296d] <= 8'he5;
		memory[16'h296e] <= 8'h51;
		memory[16'h296f] <= 8'hd8;
		memory[16'h2970] <= 8'h74;
		memory[16'h2971] <= 8'h60;
		memory[16'h2972] <= 8'h6d;
		memory[16'h2973] <= 8'h5c;
		memory[16'h2974] <= 8'hfc;
		memory[16'h2975] <= 8'h4f;
		memory[16'h2976] <= 8'hc7;
		memory[16'h2977] <= 8'h31;
		memory[16'h2978] <= 8'h18;
		memory[16'h2979] <= 8'hfc;
		memory[16'h297a] <= 8'h94;
		memory[16'h297b] <= 8'h92;
		memory[16'h297c] <= 8'ha4;
		memory[16'h297d] <= 8'hab;
		memory[16'h297e] <= 8'h90;
		memory[16'h297f] <= 8'hab;
		memory[16'h2980] <= 8'hfd;
		memory[16'h2981] <= 8'hff;
		memory[16'h2982] <= 8'h95;
		memory[16'h2983] <= 8'h73;
		memory[16'h2984] <= 8'hfd;
		memory[16'h2985] <= 8'hdb;
		memory[16'h2986] <= 8'h24;
		memory[16'h2987] <= 8'h9f;
		memory[16'h2988] <= 8'hee;
		memory[16'h2989] <= 8'hf2;
		memory[16'h298a] <= 8'h38;
		memory[16'h298b] <= 8'haa;
		memory[16'h298c] <= 8'hd7;
		memory[16'h298d] <= 8'h8a;
		memory[16'h298e] <= 8'h82;
		memory[16'h298f] <= 8'h4b;
		memory[16'h2990] <= 8'hea;
		memory[16'h2991] <= 8'hef;
		memory[16'h2992] <= 8'ha8;
		memory[16'h2993] <= 8'he7;
		memory[16'h2994] <= 8'h3f;
		memory[16'h2995] <= 8'h6f;
		memory[16'h2996] <= 8'h18;
		memory[16'h2997] <= 8'h57;
		memory[16'h2998] <= 8'h6b;
		memory[16'h2999] <= 8'had;
		memory[16'h299a] <= 8'hea;
		memory[16'h299b] <= 8'hf;
		memory[16'h299c] <= 8'h58;
		memory[16'h299d] <= 8'h7a;
		memory[16'h299e] <= 8'hbb;
		memory[16'h299f] <= 8'h55;
		memory[16'h29a0] <= 8'h79;
		memory[16'h29a1] <= 8'h50;
		memory[16'h29a2] <= 8'hc9;
		memory[16'h29a3] <= 8'h76;
		memory[16'h29a4] <= 8'h2b;
		memory[16'h29a5] <= 8'hed;
		memory[16'h29a6] <= 8'h15;
		memory[16'h29a7] <= 8'h19;
		memory[16'h29a8] <= 8'hdf;
		memory[16'h29a9] <= 8'h4e;
		memory[16'h29aa] <= 8'hc3;
		memory[16'h29ab] <= 8'hb6;
		memory[16'h29ac] <= 8'hd8;
		memory[16'h29ad] <= 8'h46;
		memory[16'h29ae] <= 8'h2;
		memory[16'h29af] <= 8'hc2;
		memory[16'h29b0] <= 8'h35;
		memory[16'h29b1] <= 8'haa;
		memory[16'h29b2] <= 8'ha9;
		memory[16'h29b3] <= 8'h74;
		memory[16'h29b4] <= 8'h19;
		memory[16'h29b5] <= 8'hc2;
		memory[16'h29b6] <= 8'hcc;
		memory[16'h29b7] <= 8'h84;
		memory[16'h29b8] <= 8'h6f;
		memory[16'h29b9] <= 8'hb6;
		memory[16'h29ba] <= 8'h93;
		memory[16'h29bb] <= 8'hc7;
		memory[16'h29bc] <= 8'h30;
		memory[16'h29bd] <= 8'h4e;
		memory[16'h29be] <= 8'h1c;
		memory[16'h29bf] <= 8'ha9;
		memory[16'h29c0] <= 8'h9f;
		memory[16'h29c1] <= 8'he5;
		memory[16'h29c2] <= 8'h1f;
		memory[16'h29c3] <= 8'hca;
		memory[16'h29c4] <= 8'hd3;
		memory[16'h29c5] <= 8'h35;
		memory[16'h29c6] <= 8'he4;
		memory[16'h29c7] <= 8'hb2;
		memory[16'h29c8] <= 8'h83;
		memory[16'h29c9] <= 8'ha7;
		memory[16'h29ca] <= 8'h69;
		memory[16'h29cb] <= 8'h5b;
		memory[16'h29cc] <= 8'hed;
		memory[16'h29cd] <= 8'h6b;
		memory[16'h29ce] <= 8'h1d;
		memory[16'h29cf] <= 8'h23;
		memory[16'h29d0] <= 8'h15;
		memory[16'h29d1] <= 8'hc7;
		memory[16'h29d2] <= 8'h97;
		memory[16'h29d3] <= 8'h2e;
		memory[16'h29d4] <= 8'h89;
		memory[16'h29d5] <= 8'h63;
		memory[16'h29d6] <= 8'hb2;
		memory[16'h29d7] <= 8'hf8;
		memory[16'h29d8] <= 8'h19;
		memory[16'h29d9] <= 8'h45;
		memory[16'h29da] <= 8'hbf;
		memory[16'h29db] <= 8'h49;
		memory[16'h29dc] <= 8'h94;
		memory[16'h29dd] <= 8'hdb;
		memory[16'h29de] <= 8'hf2;
		memory[16'h29df] <= 8'h33;
		memory[16'h29e0] <= 8'hc1;
		memory[16'h29e1] <= 8'h12;
		memory[16'h29e2] <= 8'hfd;
		memory[16'h29e3] <= 8'h94;
		memory[16'h29e4] <= 8'h47;
		memory[16'h29e5] <= 8'he1;
		memory[16'h29e6] <= 8'h46;
		memory[16'h29e7] <= 8'hca;
		memory[16'h29e8] <= 8'h89;
		memory[16'h29e9] <= 8'haf;
		memory[16'h29ea] <= 8'h25;
		memory[16'h29eb] <= 8'h76;
		memory[16'h29ec] <= 8'h1a;
		memory[16'h29ed] <= 8'h42;
		memory[16'h29ee] <= 8'h99;
		memory[16'h29ef] <= 8'h2f;
		memory[16'h29f0] <= 8'h9;
		memory[16'h29f1] <= 8'h31;
		memory[16'h29f2] <= 8'h5d;
		memory[16'h29f3] <= 8'h92;
		memory[16'h29f4] <= 8'h94;
		memory[16'h29f5] <= 8'hf;
		memory[16'h29f6] <= 8'h8a;
		memory[16'h29f7] <= 8'hae;
		memory[16'h29f8] <= 8'h55;
		memory[16'h29f9] <= 8'h49;
		memory[16'h29fa] <= 8'hf7;
		memory[16'h29fb] <= 8'he9;
		memory[16'h29fc] <= 8'h25;
		memory[16'h29fd] <= 8'hea;
		memory[16'h29fe] <= 8'h1c;
		memory[16'h29ff] <= 8'he6;
		memory[16'h2a00] <= 8'hfc;
		memory[16'h2a01] <= 8'h19;
		memory[16'h2a02] <= 8'h7a;
		memory[16'h2a03] <= 8'h43;
		memory[16'h2a04] <= 8'hfb;
		memory[16'h2a05] <= 8'hc0;
		memory[16'h2a06] <= 8'hd;
		memory[16'h2a07] <= 8'h84;
		memory[16'h2a08] <= 8'h70;
		memory[16'h2a09] <= 8'h32;
		memory[16'h2a0a] <= 8'hfa;
		memory[16'h2a0b] <= 8'h8a;
		memory[16'h2a0c] <= 8'h74;
		memory[16'h2a0d] <= 8'h94;
		memory[16'h2a0e] <= 8'hba;
		memory[16'h2a0f] <= 8'h7e;
		memory[16'h2a10] <= 8'hc5;
		memory[16'h2a11] <= 8'h17;
		memory[16'h2a12] <= 8'h10;
		memory[16'h2a13] <= 8'h59;
		memory[16'h2a14] <= 8'h27;
		memory[16'h2a15] <= 8'h9b;
		memory[16'h2a16] <= 8'h7;
		memory[16'h2a17] <= 8'h7c;
		memory[16'h2a18] <= 8'he4;
		memory[16'h2a19] <= 8'hff;
		memory[16'h2a1a] <= 8'h65;
		memory[16'h2a1b] <= 8'h9;
		memory[16'h2a1c] <= 8'he9;
		memory[16'h2a1d] <= 8'h81;
		memory[16'h2a1e] <= 8'hef;
		memory[16'h2a1f] <= 8'he5;
		memory[16'h2a20] <= 8'h9a;
		memory[16'h2a21] <= 8'h69;
		memory[16'h2a22] <= 8'h28;
		memory[16'h2a23] <= 8'h95;
		memory[16'h2a24] <= 8'h2a;
		memory[16'h2a25] <= 8'h35;
		memory[16'h2a26] <= 8'h19;
		memory[16'h2a27] <= 8'h9a;
		memory[16'h2a28] <= 8'h67;
		memory[16'h2a29] <= 8'h14;
		memory[16'h2a2a] <= 8'h24;
		memory[16'h2a2b] <= 8'hdb;
		memory[16'h2a2c] <= 8'ha8;
		memory[16'h2a2d] <= 8'hde;
		memory[16'h2a2e] <= 8'h59;
		memory[16'h2a2f] <= 8'h6d;
		memory[16'h2a30] <= 8'hf6;
		memory[16'h2a31] <= 8'h6a;
		memory[16'h2a32] <= 8'hc6;
		memory[16'h2a33] <= 8'h1d;
		memory[16'h2a34] <= 8'h5;
		memory[16'h2a35] <= 8'hce;
		memory[16'h2a36] <= 8'h99;
		memory[16'h2a37] <= 8'he9;
		memory[16'h2a38] <= 8'hcd;
		memory[16'h2a39] <= 8'hfe;
		memory[16'h2a3a] <= 8'hf3;
		memory[16'h2a3b] <= 8'hb6;
		memory[16'h2a3c] <= 8'h7f;
		memory[16'h2a3d] <= 8'he2;
		memory[16'h2a3e] <= 8'h9b;
		memory[16'h2a3f] <= 8'h19;
		memory[16'h2a40] <= 8'h4c;
		memory[16'h2a41] <= 8'hc3;
		memory[16'h2a42] <= 8'haf;
		memory[16'h2a43] <= 8'h76;
		memory[16'h2a44] <= 8'hf8;
		memory[16'h2a45] <= 8'hc8;
		memory[16'h2a46] <= 8'h10;
		memory[16'h2a47] <= 8'h5f;
		memory[16'h2a48] <= 8'hdc;
		memory[16'h2a49] <= 8'h34;
		memory[16'h2a4a] <= 8'h3a;
		memory[16'h2a4b] <= 8'h84;
		memory[16'h2a4c] <= 8'h13;
		memory[16'h2a4d] <= 8'h94;
		memory[16'h2a4e] <= 8'hf1;
		memory[16'h2a4f] <= 8'h9;
		memory[16'h2a50] <= 8'hfe;
		memory[16'h2a51] <= 8'hb8;
		memory[16'h2a52] <= 8'h26;
		memory[16'h2a53] <= 8'h3;
		memory[16'h2a54] <= 8'h86;
		memory[16'h2a55] <= 8'hbf;
		memory[16'h2a56] <= 8'hec;
		memory[16'h2a57] <= 8'h53;
		memory[16'h2a58] <= 8'hbd;
		memory[16'h2a59] <= 8'hdf;
		memory[16'h2a5a] <= 8'h9;
		memory[16'h2a5b] <= 8'h3c;
		memory[16'h2a5c] <= 8'hc2;
		memory[16'h2a5d] <= 8'ha4;
		memory[16'h2a5e] <= 8'h55;
		memory[16'h2a5f] <= 8'he;
		memory[16'h2a60] <= 8'h67;
		memory[16'h2a61] <= 8'h4;
		memory[16'h2a62] <= 8'h84;
		memory[16'h2a63] <= 8'h5f;
		memory[16'h2a64] <= 8'hcd;
		memory[16'h2a65] <= 8'h94;
		memory[16'h2a66] <= 8'hbe;
		memory[16'h2a67] <= 8'ha9;
		memory[16'h2a68] <= 8'hc8;
		memory[16'h2a69] <= 8'hf8;
		memory[16'h2a6a] <= 8'h2e;
		memory[16'h2a6b] <= 8'hdb;
		memory[16'h2a6c] <= 8'h8c;
		memory[16'h2a6d] <= 8'h1f;
		memory[16'h2a6e] <= 8'he4;
		memory[16'h2a6f] <= 8'h8a;
		memory[16'h2a70] <= 8'hd7;
		memory[16'h2a71] <= 8'ha;
		memory[16'h2a72] <= 8'h8d;
		memory[16'h2a73] <= 8'h5d;
		memory[16'h2a74] <= 8'hc9;
		memory[16'h2a75] <= 8'h7a;
		memory[16'h2a76] <= 8'hb0;
		memory[16'h2a77] <= 8'h86;
		memory[16'h2a78] <= 8'h59;
		memory[16'h2a79] <= 8'hb9;
		memory[16'h2a7a] <= 8'hc2;
		memory[16'h2a7b] <= 8'h1b;
		memory[16'h2a7c] <= 8'h5d;
		memory[16'h2a7d] <= 8'h18;
		memory[16'h2a7e] <= 8'h29;
		memory[16'h2a7f] <= 8'hc4;
		memory[16'h2a80] <= 8'h1c;
		memory[16'h2a81] <= 8'had;
		memory[16'h2a82] <= 8'h23;
		memory[16'h2a83] <= 8'he9;
		memory[16'h2a84] <= 8'h41;
		memory[16'h2a85] <= 8'he1;
		memory[16'h2a86] <= 8'h93;
		memory[16'h2a87] <= 8'ha;
		memory[16'h2a88] <= 8'hda;
		memory[16'h2a89] <= 8'hc1;
		memory[16'h2a8a] <= 8'he5;
		memory[16'h2a8b] <= 8'h66;
		memory[16'h2a8c] <= 8'he0;
		memory[16'h2a8d] <= 8'hca;
		memory[16'h2a8e] <= 8'hf1;
		memory[16'h2a8f] <= 8'hb8;
		memory[16'h2a90] <= 8'hd4;
		memory[16'h2a91] <= 8'h7e;
		memory[16'h2a92] <= 8'h15;
		memory[16'h2a93] <= 8'h9e;
		memory[16'h2a94] <= 8'hf8;
		memory[16'h2a95] <= 8'hc6;
		memory[16'h2a96] <= 8'h24;
		memory[16'h2a97] <= 8'h52;
		memory[16'h2a98] <= 8'h7f;
		memory[16'h2a99] <= 8'he7;
		memory[16'h2a9a] <= 8'h6d;
		memory[16'h2a9b] <= 8'hdd;
		memory[16'h2a9c] <= 8'hff;
		memory[16'h2a9d] <= 8'h97;
		memory[16'h2a9e] <= 8'ha1;
		memory[16'h2a9f] <= 8'h1b;
		memory[16'h2aa0] <= 8'h44;
		memory[16'h2aa1] <= 8'hc5;
		memory[16'h2aa2] <= 8'h5;
		memory[16'h2aa3] <= 8'h86;
		memory[16'h2aa4] <= 8'ha6;
		memory[16'h2aa5] <= 8'h98;
		memory[16'h2aa6] <= 8'h90;
		memory[16'h2aa7] <= 8'h80;
		memory[16'h2aa8] <= 8'h59;
		memory[16'h2aa9] <= 8'h75;
		memory[16'h2aaa] <= 8'he7;
		memory[16'h2aab] <= 8'h39;
		memory[16'h2aac] <= 8'h3f;
		memory[16'h2aad] <= 8'hd8;
		memory[16'h2aae] <= 8'hf1;
		memory[16'h2aaf] <= 8'h14;
		memory[16'h2ab0] <= 8'h56;
		memory[16'h2ab1] <= 8'h7;
		memory[16'h2ab2] <= 8'hb2;
		memory[16'h2ab3] <= 8'h4f;
		memory[16'h2ab4] <= 8'hcd;
		memory[16'h2ab5] <= 8'hd6;
		memory[16'h2ab6] <= 8'ha1;
		memory[16'h2ab7] <= 8'h4c;
		memory[16'h2ab8] <= 8'hbd;
		memory[16'h2ab9] <= 8'he;
		memory[16'h2aba] <= 8'h29;
		memory[16'h2abb] <= 8'hbc;
		memory[16'h2abc] <= 8'ha5;
		memory[16'h2abd] <= 8'hcb;
		memory[16'h2abe] <= 8'hd8;
		memory[16'h2abf] <= 8'hea;
		memory[16'h2ac0] <= 8'h90;
		memory[16'h2ac1] <= 8'hdd;
		memory[16'h2ac2] <= 8'h70;
		memory[16'h2ac3] <= 8'h36;
		memory[16'h2ac4] <= 8'h75;
		memory[16'h2ac5] <= 8'h0;
		memory[16'h2ac6] <= 8'hb7;
		memory[16'h2ac7] <= 8'hce;
		memory[16'h2ac8] <= 8'h75;
		memory[16'h2ac9] <= 8'h9e;
		memory[16'h2aca] <= 8'h7;
		memory[16'h2acb] <= 8'hb5;
		memory[16'h2acc] <= 8'h76;
		memory[16'h2acd] <= 8'hf9;
		memory[16'h2ace] <= 8'hc9;
		memory[16'h2acf] <= 8'hcc;
		memory[16'h2ad0] <= 8'h0;
		memory[16'h2ad1] <= 8'h7b;
		memory[16'h2ad2] <= 8'h1b;
		memory[16'h2ad3] <= 8'hcd;
		memory[16'h2ad4] <= 8'h51;
		memory[16'h2ad5] <= 8'hbc;
		memory[16'h2ad6] <= 8'h19;
		memory[16'h2ad7] <= 8'hf;
		memory[16'h2ad8] <= 8'hcb;
		memory[16'h2ad9] <= 8'h43;
		memory[16'h2ada] <= 8'hcb;
		memory[16'h2adb] <= 8'h70;
		memory[16'h2adc] <= 8'he;
		memory[16'h2add] <= 8'ha3;
		memory[16'h2ade] <= 8'h5a;
		memory[16'h2adf] <= 8'h9e;
		memory[16'h2ae0] <= 8'h80;
		memory[16'h2ae1] <= 8'hca;
		memory[16'h2ae2] <= 8'hd4;
		memory[16'h2ae3] <= 8'hf5;
		memory[16'h2ae4] <= 8'hca;
		memory[16'h2ae5] <= 8'h8b;
		memory[16'h2ae6] <= 8'hc3;
		memory[16'h2ae7] <= 8'h40;
		memory[16'h2ae8] <= 8'h29;
		memory[16'h2ae9] <= 8'hcb;
		memory[16'h2aea] <= 8'hf5;
		memory[16'h2aeb] <= 8'h9f;
		memory[16'h2aec] <= 8'hc4;
		memory[16'h2aed] <= 8'hbe;
		memory[16'h2aee] <= 8'h6c;
		memory[16'h2aef] <= 8'hc4;
		memory[16'h2af0] <= 8'h39;
		memory[16'h2af1] <= 8'h87;
		memory[16'h2af2] <= 8'h91;
		memory[16'h2af3] <= 8'h8a;
		memory[16'h2af4] <= 8'h44;
		memory[16'h2af5] <= 8'haa;
		memory[16'h2af6] <= 8'h99;
		memory[16'h2af7] <= 8'hf;
		memory[16'h2af8] <= 8'hed;
		memory[16'h2af9] <= 8'h65;
		memory[16'h2afa] <= 8'h7f;
		memory[16'h2afb] <= 8'hfb;
		memory[16'h2afc] <= 8'h8;
		memory[16'h2afd] <= 8'hda;
		memory[16'h2afe] <= 8'h99;
		memory[16'h2aff] <= 8'h89;
		memory[16'h2b00] <= 8'ha4;
		memory[16'h2b01] <= 8'h6e;
		memory[16'h2b02] <= 8'h7e;
		memory[16'h2b03] <= 8'h6f;
		memory[16'h2b04] <= 8'hf9;
		memory[16'h2b05] <= 8'h42;
		memory[16'h2b06] <= 8'haf;
		memory[16'h2b07] <= 8'h23;
		memory[16'h2b08] <= 8'hd;
		memory[16'h2b09] <= 8'ha4;
		memory[16'h2b0a] <= 8'hc2;
		memory[16'h2b0b] <= 8'hd1;
		memory[16'h2b0c] <= 8'h62;
		memory[16'h2b0d] <= 8'h2e;
		memory[16'h2b0e] <= 8'h95;
		memory[16'h2b0f] <= 8'h9b;
		memory[16'h2b10] <= 8'hb6;
		memory[16'h2b11] <= 8'h26;
		memory[16'h2b12] <= 8'h25;
		memory[16'h2b13] <= 8'hfa;
		memory[16'h2b14] <= 8'hd0;
		memory[16'h2b15] <= 8'hbf;
		memory[16'h2b16] <= 8'h9;
		memory[16'h2b17] <= 8'hbe;
		memory[16'h2b18] <= 8'h24;
		memory[16'h2b19] <= 8'h88;
		memory[16'h2b1a] <= 8'hb9;
		memory[16'h2b1b] <= 8'h2c;
		memory[16'h2b1c] <= 8'h62;
		memory[16'h2b1d] <= 8'h53;
		memory[16'h2b1e] <= 8'hb5;
		memory[16'h2b1f] <= 8'h7;
		memory[16'h2b20] <= 8'hc1;
		memory[16'h2b21] <= 8'h34;
		memory[16'h2b22] <= 8'h76;
		memory[16'h2b23] <= 8'hba;
		memory[16'h2b24] <= 8'h76;
		memory[16'h2b25] <= 8'h25;
		memory[16'h2b26] <= 8'hdd;
		memory[16'h2b27] <= 8'h83;
		memory[16'h2b28] <= 8'hc9;
		memory[16'h2b29] <= 8'ha0;
		memory[16'h2b2a] <= 8'h54;
		memory[16'h2b2b] <= 8'h2b;
		memory[16'h2b2c] <= 8'hce;
		memory[16'h2b2d] <= 8'he9;
		memory[16'h2b2e] <= 8'hc6;
		memory[16'h2b2f] <= 8'h84;
		memory[16'h2b30] <= 8'hf;
		memory[16'h2b31] <= 8'heb;
		memory[16'h2b32] <= 8'h7e;
		memory[16'h2b33] <= 8'hdf;
		memory[16'h2b34] <= 8'haa;
		memory[16'h2b35] <= 8'h87;
		memory[16'h2b36] <= 8'h9d;
		memory[16'h2b37] <= 8'hce;
		memory[16'h2b38] <= 8'h10;
		memory[16'h2b39] <= 8'h57;
		memory[16'h2b3a] <= 8'hfb;
		memory[16'h2b3b] <= 8'h72;
		memory[16'h2b3c] <= 8'haa;
		memory[16'h2b3d] <= 8'hb0;
		memory[16'h2b3e] <= 8'h79;
		memory[16'h2b3f] <= 8'h6b;
		memory[16'h2b40] <= 8'he4;
		memory[16'h2b41] <= 8'hef;
		memory[16'h2b42] <= 8'h25;
		memory[16'h2b43] <= 8'h5a;
		memory[16'h2b44] <= 8'h14;
		memory[16'h2b45] <= 8'h3;
		memory[16'h2b46] <= 8'hdd;
		memory[16'h2b47] <= 8'hdd;
		memory[16'h2b48] <= 8'ha3;
		memory[16'h2b49] <= 8'h31;
		memory[16'h2b4a] <= 8'h8;
		memory[16'h2b4b] <= 8'h71;
		memory[16'h2b4c] <= 8'h1a;
		memory[16'h2b4d] <= 8'hce;
		memory[16'h2b4e] <= 8'hf6;
		memory[16'h2b4f] <= 8'h29;
		memory[16'h2b50] <= 8'hba;
		memory[16'h2b51] <= 8'h74;
		memory[16'h2b52] <= 8'h9;
		memory[16'h2b53] <= 8'h64;
		memory[16'h2b54] <= 8'hfc;
		memory[16'h2b55] <= 8'ha6;
		memory[16'h2b56] <= 8'h33;
		memory[16'h2b57] <= 8'hc;
		memory[16'h2b58] <= 8'hfd;
		memory[16'h2b59] <= 8'h2e;
		memory[16'h2b5a] <= 8'h7e;
		memory[16'h2b5b] <= 8'ha7;
		memory[16'h2b5c] <= 8'hde;
		memory[16'h2b5d] <= 8'hf8;
		memory[16'h2b5e] <= 8'h12;
		memory[16'h2b5f] <= 8'hc3;
		memory[16'h2b60] <= 8'he7;
		memory[16'h2b61] <= 8'h38;
		memory[16'h2b62] <= 8'h1d;
		memory[16'h2b63] <= 8'hfc;
		memory[16'h2b64] <= 8'h3b;
		memory[16'h2b65] <= 8'hfb;
		memory[16'h2b66] <= 8'hd9;
		memory[16'h2b67] <= 8'hde;
		memory[16'h2b68] <= 8'h2c;
		memory[16'h2b69] <= 8'he2;
		memory[16'h2b6a] <= 8'h4f;
		memory[16'h2b6b] <= 8'h47;
		memory[16'h2b6c] <= 8'hb0;
		memory[16'h2b6d] <= 8'h45;
		memory[16'h2b6e] <= 8'h70;
		memory[16'h2b6f] <= 8'h6a;
		memory[16'h2b70] <= 8'hba;
		memory[16'h2b71] <= 8'h79;
		memory[16'h2b72] <= 8'hcf;
		memory[16'h2b73] <= 8'hb6;
		memory[16'h2b74] <= 8'h20;
		memory[16'h2b75] <= 8'h2;
		memory[16'h2b76] <= 8'hc2;
		memory[16'h2b77] <= 8'h1d;
		memory[16'h2b78] <= 8'h30;
		memory[16'h2b79] <= 8'h40;
		memory[16'h2b7a] <= 8'hc5;
		memory[16'h2b7b] <= 8'he;
		memory[16'h2b7c] <= 8'h38;
		memory[16'h2b7d] <= 8'hd7;
		memory[16'h2b7e] <= 8'hd1;
		memory[16'h2b7f] <= 8'h20;
		memory[16'h2b80] <= 8'hf;
		memory[16'h2b81] <= 8'hef;
		memory[16'h2b82] <= 8'h1c;
		memory[16'h2b83] <= 8'h4a;
		memory[16'h2b84] <= 8'hea;
		memory[16'h2b85] <= 8'hf5;
		memory[16'h2b86] <= 8'h28;
		memory[16'h2b87] <= 8'h16;
		memory[16'h2b88] <= 8'hd7;
		memory[16'h2b89] <= 8'h78;
		memory[16'h2b8a] <= 8'h5d;
		memory[16'h2b8b] <= 8'h88;
		memory[16'h2b8c] <= 8'hbd;
		memory[16'h2b8d] <= 8'hce;
		memory[16'h2b8e] <= 8'hf2;
		memory[16'h2b8f] <= 8'h77;
		memory[16'h2b90] <= 8'h47;
		memory[16'h2b91] <= 8'hc1;
		memory[16'h2b92] <= 8'h2d;
		memory[16'h2b93] <= 8'h67;
		memory[16'h2b94] <= 8'hc3;
		memory[16'h2b95] <= 8'hef;
		memory[16'h2b96] <= 8'h85;
		memory[16'h2b97] <= 8'hf3;
		memory[16'h2b98] <= 8'h30;
		memory[16'h2b99] <= 8'h4a;
		memory[16'h2b9a] <= 8'h2;
		memory[16'h2b9b] <= 8'h68;
		memory[16'h2b9c] <= 8'h21;
		memory[16'h2b9d] <= 8'hd3;
		memory[16'h2b9e] <= 8'h88;
		memory[16'h2b9f] <= 8'h31;
		memory[16'h2ba0] <= 8'hc2;
		memory[16'h2ba1] <= 8'ha4;
		memory[16'h2ba2] <= 8'h7b;
		memory[16'h2ba3] <= 8'hac;
		memory[16'h2ba4] <= 8'h9a;
		memory[16'h2ba5] <= 8'ha4;
		memory[16'h2ba6] <= 8'hc3;
		memory[16'h2ba7] <= 8'h71;
		memory[16'h2ba8] <= 8'h1c;
		memory[16'h2ba9] <= 8'h20;
		memory[16'h2baa] <= 8'hf9;
		memory[16'h2bab] <= 8'hd9;
		memory[16'h2bac] <= 8'hee;
		memory[16'h2bad] <= 8'hec;
		memory[16'h2bae] <= 8'h51;
		memory[16'h2baf] <= 8'h36;
		memory[16'h2bb0] <= 8'had;
		memory[16'h2bb1] <= 8'h7e;
		memory[16'h2bb2] <= 8'h9d;
		memory[16'h2bb3] <= 8'h71;
		memory[16'h2bb4] <= 8'h6e;
		memory[16'h2bb5] <= 8'h22;
		memory[16'h2bb6] <= 8'h64;
		memory[16'h2bb7] <= 8'h9e;
		memory[16'h2bb8] <= 8'h6c;
		memory[16'h2bb9] <= 8'h66;
		memory[16'h2bba] <= 8'h6;
		memory[16'h2bbb] <= 8'h8e;
		memory[16'h2bbc] <= 8'h3a;
		memory[16'h2bbd] <= 8'h8f;
		memory[16'h2bbe] <= 8'hbf;
		memory[16'h2bbf] <= 8'hfc;
		memory[16'h2bc0] <= 8'h33;
		memory[16'h2bc1] <= 8'h3a;
		memory[16'h2bc2] <= 8'ha9;
		memory[16'h2bc3] <= 8'hcd;
		memory[16'h2bc4] <= 8'hde;
		memory[16'h2bc5] <= 8'h6c;
		memory[16'h2bc6] <= 8'h3f;
		memory[16'h2bc7] <= 8'hfa;
		memory[16'h2bc8] <= 8'h8c;
		memory[16'h2bc9] <= 8'h38;
		memory[16'h2bca] <= 8'hd4;
		memory[16'h2bcb] <= 8'h7b;
		memory[16'h2bcc] <= 8'h24;
		memory[16'h2bcd] <= 8'h25;
		memory[16'h2bce] <= 8'hb1;
		memory[16'h2bcf] <= 8'hd2;
		memory[16'h2bd0] <= 8'ha3;
		memory[16'h2bd1] <= 8'h4e;
		memory[16'h2bd2] <= 8'h43;
		memory[16'h2bd3] <= 8'h11;
		memory[16'h2bd4] <= 8'h71;
		memory[16'h2bd5] <= 8'ha7;
		memory[16'h2bd6] <= 8'haf;
		memory[16'h2bd7] <= 8'hdd;
		memory[16'h2bd8] <= 8'he;
		memory[16'h2bd9] <= 8'hb6;
		memory[16'h2bda] <= 8'h6b;
		memory[16'h2bdb] <= 8'h48;
		memory[16'h2bdc] <= 8'h45;
		memory[16'h2bdd] <= 8'h2a;
		memory[16'h2bde] <= 8'h44;
		memory[16'h2bdf] <= 8'h78;
		memory[16'h2be0] <= 8'h65;
		memory[16'h2be1] <= 8'hed;
		memory[16'h2be2] <= 8'h46;
		memory[16'h2be3] <= 8'h43;
		memory[16'h2be4] <= 8'h59;
		memory[16'h2be5] <= 8'h85;
		memory[16'h2be6] <= 8'h3e;
		memory[16'h2be7] <= 8'he6;
		memory[16'h2be8] <= 8'hbd;
		memory[16'h2be9] <= 8'h12;
		memory[16'h2bea] <= 8'h61;
		memory[16'h2beb] <= 8'he2;
		memory[16'h2bec] <= 8'h37;
		memory[16'h2bed] <= 8'h12;
		memory[16'h2bee] <= 8'hb4;
		memory[16'h2bef] <= 8'hda;
		memory[16'h2bf0] <= 8'h60;
		memory[16'h2bf1] <= 8'hf7;
		memory[16'h2bf2] <= 8'hec;
		memory[16'h2bf3] <= 8'hd1;
		memory[16'h2bf4] <= 8'h9e;
		memory[16'h2bf5] <= 8'h9b;
		memory[16'h2bf6] <= 8'haf;
		memory[16'h2bf7] <= 8'hac;
		memory[16'h2bf8] <= 8'h51;
		memory[16'h2bf9] <= 8'h1a;
		memory[16'h2bfa] <= 8'hf4;
		memory[16'h2bfb] <= 8'h96;
		memory[16'h2bfc] <= 8'h45;
		memory[16'h2bfd] <= 8'h39;
		memory[16'h2bfe] <= 8'hf;
		memory[16'h2bff] <= 8'haa;
		memory[16'h2c00] <= 8'h26;
		memory[16'h2c01] <= 8'h55;
		memory[16'h2c02] <= 8'hed;
		memory[16'h2c03] <= 8'h80;
		memory[16'h2c04] <= 8'hda;
		memory[16'h2c05] <= 8'h2b;
		memory[16'h2c06] <= 8'h66;
		memory[16'h2c07] <= 8'h97;
		memory[16'h2c08] <= 8'h3d;
		memory[16'h2c09] <= 8'hc7;
		memory[16'h2c0a] <= 8'h79;
		memory[16'h2c0b] <= 8'h74;
		memory[16'h2c0c] <= 8'hd9;
		memory[16'h2c0d] <= 8'h2d;
		memory[16'h2c0e] <= 8'h4f;
		memory[16'h2c0f] <= 8'h39;
		memory[16'h2c10] <= 8'h24;
		memory[16'h2c11] <= 8'h3b;
		memory[16'h2c12] <= 8'hb;
		memory[16'h2c13] <= 8'hc3;
		memory[16'h2c14] <= 8'hd6;
		memory[16'h2c15] <= 8'hba;
		memory[16'h2c16] <= 8'h6f;
		memory[16'h2c17] <= 8'h28;
		memory[16'h2c18] <= 8'hd4;
		memory[16'h2c19] <= 8'h64;
		memory[16'h2c1a] <= 8'hbe;
		memory[16'h2c1b] <= 8'h19;
		memory[16'h2c1c] <= 8'h9d;
		memory[16'h2c1d] <= 8'hcd;
		memory[16'h2c1e] <= 8'hc3;
		memory[16'h2c1f] <= 8'hc3;
		memory[16'h2c20] <= 8'h22;
		memory[16'h2c21] <= 8'hb1;
		memory[16'h2c22] <= 8'h43;
		memory[16'h2c23] <= 8'hfc;
		memory[16'h2c24] <= 8'hdc;
		memory[16'h2c25] <= 8'ha9;
		memory[16'h2c26] <= 8'h94;
		memory[16'h2c27] <= 8'h1a;
		memory[16'h2c28] <= 8'h70;
		memory[16'h2c29] <= 8'hd;
		memory[16'h2c2a] <= 8'h8e;
		memory[16'h2c2b] <= 8'h49;
		memory[16'h2c2c] <= 8'h3b;
		memory[16'h2c2d] <= 8'hdd;
		memory[16'h2c2e] <= 8'h83;
		memory[16'h2c2f] <= 8'h5f;
		memory[16'h2c30] <= 8'h18;
		memory[16'h2c31] <= 8'h8e;
		memory[16'h2c32] <= 8'h22;
		memory[16'h2c33] <= 8'hef;
		memory[16'h2c34] <= 8'h48;
		memory[16'h2c35] <= 8'h92;
		memory[16'h2c36] <= 8'h17;
		memory[16'h2c37] <= 8'h1c;
		memory[16'h2c38] <= 8'hf6;
		memory[16'h2c39] <= 8'hd5;
		memory[16'h2c3a] <= 8'h36;
		memory[16'h2c3b] <= 8'h93;
		memory[16'h2c3c] <= 8'ha3;
		memory[16'h2c3d] <= 8'hf9;
		memory[16'h2c3e] <= 8'h56;
		memory[16'h2c3f] <= 8'hc5;
		memory[16'h2c40] <= 8'haa;
		memory[16'h2c41] <= 8'h9a;
		memory[16'h2c42] <= 8'hc2;
		memory[16'h2c43] <= 8'h87;
		memory[16'h2c44] <= 8'h43;
		memory[16'h2c45] <= 8'h56;
		memory[16'h2c46] <= 8'ha1;
		memory[16'h2c47] <= 8'hb4;
		memory[16'h2c48] <= 8'h63;
		memory[16'h2c49] <= 8'h2f;
		memory[16'h2c4a] <= 8'hfd;
		memory[16'h2c4b] <= 8'h9e;
		memory[16'h2c4c] <= 8'hd;
		memory[16'h2c4d] <= 8'h80;
		memory[16'h2c4e] <= 8'hfe;
		memory[16'h2c4f] <= 8'h25;
		memory[16'h2c50] <= 8'he;
		memory[16'h2c51] <= 8'h20;
		memory[16'h2c52] <= 8'h14;
		memory[16'h2c53] <= 8'h56;
		memory[16'h2c54] <= 8'hb2;
		memory[16'h2c55] <= 8'h2b;
		memory[16'h2c56] <= 8'h73;
		memory[16'h2c57] <= 8'ha8;
		memory[16'h2c58] <= 8'h1;
		memory[16'h2c59] <= 8'ha9;
		memory[16'h2c5a] <= 8'h3b;
		memory[16'h2c5b] <= 8'ha4;
		memory[16'h2c5c] <= 8'ha2;
		memory[16'h2c5d] <= 8'h92;
		memory[16'h2c5e] <= 8'h69;
		memory[16'h2c5f] <= 8'h4d;
		memory[16'h2c60] <= 8'h2c;
		memory[16'h2c61] <= 8'h2b;
		memory[16'h2c62] <= 8'hd4;
		memory[16'h2c63] <= 8'h6f;
		memory[16'h2c64] <= 8'h81;
		memory[16'h2c65] <= 8'h75;
		memory[16'h2c66] <= 8'h23;
		memory[16'h2c67] <= 8'he5;
		memory[16'h2c68] <= 8'ha4;
		memory[16'h2c69] <= 8'h21;
		memory[16'h2c6a] <= 8'h83;
		memory[16'h2c6b] <= 8'hb1;
		memory[16'h2c6c] <= 8'ha1;
		memory[16'h2c6d] <= 8'h81;
		memory[16'h2c6e] <= 8'hd7;
		memory[16'h2c6f] <= 8'hb0;
		memory[16'h2c70] <= 8'ha2;
		memory[16'h2c71] <= 8'heb;
		memory[16'h2c72] <= 8'h6;
		memory[16'h2c73] <= 8'h54;
		memory[16'h2c74] <= 8'h17;
		memory[16'h2c75] <= 8'h79;
		memory[16'h2c76] <= 8'hfd;
		memory[16'h2c77] <= 8'h18;
		memory[16'h2c78] <= 8'h22;
		memory[16'h2c79] <= 8'h38;
		memory[16'h2c7a] <= 8'hbc;
		memory[16'h2c7b] <= 8'hc5;
		memory[16'h2c7c] <= 8'hca;
		memory[16'h2c7d] <= 8'h25;
		memory[16'h2c7e] <= 8'h12;
		memory[16'h2c7f] <= 8'hf6;
		memory[16'h2c80] <= 8'h51;
		memory[16'h2c81] <= 8'he6;
		memory[16'h2c82] <= 8'h66;
		memory[16'h2c83] <= 8'hd2;
		memory[16'h2c84] <= 8'h5b;
		memory[16'h2c85] <= 8'h89;
		memory[16'h2c86] <= 8'hb7;
		memory[16'h2c87] <= 8'hff;
		memory[16'h2c88] <= 8'haa;
		memory[16'h2c89] <= 8'h3b;
		memory[16'h2c8a] <= 8'hb1;
		memory[16'h2c8b] <= 8'h4c;
		memory[16'h2c8c] <= 8'hbc;
		memory[16'h2c8d] <= 8'h88;
		memory[16'h2c8e] <= 8'hfc;
		memory[16'h2c8f] <= 8'h5e;
		memory[16'h2c90] <= 8'h73;
		memory[16'h2c91] <= 8'h2;
		memory[16'h2c92] <= 8'hb3;
		memory[16'h2c93] <= 8'h8a;
		memory[16'h2c94] <= 8'h7c;
		memory[16'h2c95] <= 8'hb0;
		memory[16'h2c96] <= 8'ha2;
		memory[16'h2c97] <= 8'h9e;
		memory[16'h2c98] <= 8'he8;
		memory[16'h2c99] <= 8'h5e;
		memory[16'h2c9a] <= 8'h63;
		memory[16'h2c9b] <= 8'hb3;
		memory[16'h2c9c] <= 8'h84;
		memory[16'h2c9d] <= 8'h75;
		memory[16'h2c9e] <= 8'ha9;
		memory[16'h2c9f] <= 8'hd5;
		memory[16'h2ca0] <= 8'h5b;
		memory[16'h2ca1] <= 8'hf;
		memory[16'h2ca2] <= 8'ha7;
		memory[16'h2ca3] <= 8'hb6;
		memory[16'h2ca4] <= 8'h99;
		memory[16'h2ca5] <= 8'h5f;
		memory[16'h2ca6] <= 8'hb6;
		memory[16'h2ca7] <= 8'h43;
		memory[16'h2ca8] <= 8'h9a;
		memory[16'h2ca9] <= 8'h67;
		memory[16'h2caa] <= 8'h8f;
		memory[16'h2cab] <= 8'h56;
		memory[16'h2cac] <= 8'hef;
		memory[16'h2cad] <= 8'h8b;
		memory[16'h2cae] <= 8'hb5;
		memory[16'h2caf] <= 8'h62;
		memory[16'h2cb0] <= 8'h8e;
		memory[16'h2cb1] <= 8'h68;
		memory[16'h2cb2] <= 8'hed;
		memory[16'h2cb3] <= 8'ha;
		memory[16'h2cb4] <= 8'h18;
		memory[16'h2cb5] <= 8'h8f;
		memory[16'h2cb6] <= 8'ha8;
		memory[16'h2cb7] <= 8'h0;
		memory[16'h2cb8] <= 8'hee;
		memory[16'h2cb9] <= 8'hc;
		memory[16'h2cba] <= 8'hb3;
		memory[16'h2cbb] <= 8'h72;
		memory[16'h2cbc] <= 8'h81;
		memory[16'h2cbd] <= 8'h5d;
		memory[16'h2cbe] <= 8'h47;
		memory[16'h2cbf] <= 8'hdd;
		memory[16'h2cc0] <= 8'h6c;
		memory[16'h2cc1] <= 8'hee;
		memory[16'h2cc2] <= 8'h93;
		memory[16'h2cc3] <= 8'h5;
		memory[16'h2cc4] <= 8'h4d;
		memory[16'h2cc5] <= 8'h49;
		memory[16'h2cc6] <= 8'h49;
		memory[16'h2cc7] <= 8'he7;
		memory[16'h2cc8] <= 8'hb0;
		memory[16'h2cc9] <= 8'hd8;
		memory[16'h2cca] <= 8'h3e;
		memory[16'h2ccb] <= 8'h9f;
		memory[16'h2ccc] <= 8'h64;
		memory[16'h2ccd] <= 8'hf3;
		memory[16'h2cce] <= 8'h2;
		memory[16'h2ccf] <= 8'hf2;
		memory[16'h2cd0] <= 8'h5b;
		memory[16'h2cd1] <= 8'hef;
		memory[16'h2cd2] <= 8'hfc;
		memory[16'h2cd3] <= 8'h73;
		memory[16'h2cd4] <= 8'h7e;
		memory[16'h2cd5] <= 8'ha4;
		memory[16'h2cd6] <= 8'h73;
		memory[16'h2cd7] <= 8'h6c;
		memory[16'h2cd8] <= 8'hb0;
		memory[16'h2cd9] <= 8'h27;
		memory[16'h2cda] <= 8'hde;
		memory[16'h2cdb] <= 8'h32;
		memory[16'h2cdc] <= 8'h84;
		memory[16'h2cdd] <= 8'h25;
		memory[16'h2cde] <= 8'hf;
		memory[16'h2cdf] <= 8'hf0;
		memory[16'h2ce0] <= 8'h14;
		memory[16'h2ce1] <= 8'ha2;
		memory[16'h2ce2] <= 8'hf6;
		memory[16'h2ce3] <= 8'h61;
		memory[16'h2ce4] <= 8'hec;
		memory[16'h2ce5] <= 8'h3f;
		memory[16'h2ce6] <= 8'h49;
		memory[16'h2ce7] <= 8'h9c;
		memory[16'h2ce8] <= 8'h17;
		memory[16'h2ce9] <= 8'h87;
		memory[16'h2cea] <= 8'h3c;
		memory[16'h2ceb] <= 8'h7b;
		memory[16'h2cec] <= 8'h7a;
		memory[16'h2ced] <= 8'h3e;
		memory[16'h2cee] <= 8'h6d;
		memory[16'h2cef] <= 8'hd5;
		memory[16'h2cf0] <= 8'h2d;
		memory[16'h2cf1] <= 8'h69;
		memory[16'h2cf2] <= 8'h48;
		memory[16'h2cf3] <= 8'hab;
		memory[16'h2cf4] <= 8'he;
		memory[16'h2cf5] <= 8'hbb;
		memory[16'h2cf6] <= 8'h18;
		memory[16'h2cf7] <= 8'hbe;
		memory[16'h2cf8] <= 8'he2;
		memory[16'h2cf9] <= 8'hf6;
		memory[16'h2cfa] <= 8'hf0;
		memory[16'h2cfb] <= 8'h66;
		memory[16'h2cfc] <= 8'h1c;
		memory[16'h2cfd] <= 8'hff;
		memory[16'h2cfe] <= 8'h57;
		memory[16'h2cff] <= 8'h30;
		memory[16'h2d00] <= 8'ha2;
		memory[16'h2d01] <= 8'h4d;
		memory[16'h2d02] <= 8'h91;
		memory[16'h2d03] <= 8'h8e;
		memory[16'h2d04] <= 8'h8c;
		memory[16'h2d05] <= 8'hda;
		memory[16'h2d06] <= 8'h2a;
		memory[16'h2d07] <= 8'ha3;
		memory[16'h2d08] <= 8'h61;
		memory[16'h2d09] <= 8'h66;
		memory[16'h2d0a] <= 8'h1f;
		memory[16'h2d0b] <= 8'hdb;
		memory[16'h2d0c] <= 8'ha4;
		memory[16'h2d0d] <= 8'h8c;
		memory[16'h2d0e] <= 8'hb0;
		memory[16'h2d0f] <= 8'hd1;
		memory[16'h2d10] <= 8'hf6;
		memory[16'h2d11] <= 8'hf8;
		memory[16'h2d12] <= 8'h7d;
		memory[16'h2d13] <= 8'h4;
		memory[16'h2d14] <= 8'hb4;
		memory[16'h2d15] <= 8'h95;
		memory[16'h2d16] <= 8'hc2;
		memory[16'h2d17] <= 8'h96;
		memory[16'h2d18] <= 8'h8b;
		memory[16'h2d19] <= 8'hb3;
		memory[16'h2d1a] <= 8'hfd;
		memory[16'h2d1b] <= 8'ha7;
		memory[16'h2d1c] <= 8'hb2;
		memory[16'h2d1d] <= 8'h54;
		memory[16'h2d1e] <= 8'hd7;
		memory[16'h2d1f] <= 8'h54;
		memory[16'h2d20] <= 8'ha1;
		memory[16'h2d21] <= 8'h69;
		memory[16'h2d22] <= 8'he2;
		memory[16'h2d23] <= 8'h2d;
		memory[16'h2d24] <= 8'h43;
		memory[16'h2d25] <= 8'hd;
		memory[16'h2d26] <= 8'hd0;
		memory[16'h2d27] <= 8'ha5;
		memory[16'h2d28] <= 8'h73;
		memory[16'h2d29] <= 8'hef;
		memory[16'h2d2a] <= 8'h80;
		memory[16'h2d2b] <= 8'h18;
		memory[16'h2d2c] <= 8'h7c;
		memory[16'h2d2d] <= 8'h31;
		memory[16'h2d2e] <= 8'he9;
		memory[16'h2d2f] <= 8'h72;
		memory[16'h2d30] <= 8'h29;
		memory[16'h2d31] <= 8'h66;
		memory[16'h2d32] <= 8'h76;
		memory[16'h2d33] <= 8'hdd;
		memory[16'h2d34] <= 8'hfb;
		memory[16'h2d35] <= 8'h38;
		memory[16'h2d36] <= 8'h74;
		memory[16'h2d37] <= 8'h87;
		memory[16'h2d38] <= 8'heb;
		memory[16'h2d39] <= 8'h71;
		memory[16'h2d3a] <= 8'h2e;
		memory[16'h2d3b] <= 8'h9e;
		memory[16'h2d3c] <= 8'hc5;
		memory[16'h2d3d] <= 8'h6;
		memory[16'h2d3e] <= 8'hf2;
		memory[16'h2d3f] <= 8'h66;
		memory[16'h2d40] <= 8'h6f;
		memory[16'h2d41] <= 8'hd5;
		memory[16'h2d42] <= 8'h93;
		memory[16'h2d43] <= 8'hb2;
		memory[16'h2d44] <= 8'he2;
		memory[16'h2d45] <= 8'h63;
		memory[16'h2d46] <= 8'h57;
		memory[16'h2d47] <= 8'h55;
		memory[16'h2d48] <= 8'h53;
		memory[16'h2d49] <= 8'hd8;
		memory[16'h2d4a] <= 8'h6d;
		memory[16'h2d4b] <= 8'hcf;
		memory[16'h2d4c] <= 8'h9;
		memory[16'h2d4d] <= 8'h57;
		memory[16'h2d4e] <= 8'h41;
		memory[16'h2d4f] <= 8'h32;
		memory[16'h2d50] <= 8'hbd;
		memory[16'h2d51] <= 8'hb7;
		memory[16'h2d52] <= 8'h10;
		memory[16'h2d53] <= 8'hb9;
		memory[16'h2d54] <= 8'hef;
		memory[16'h2d55] <= 8'h84;
		memory[16'h2d56] <= 8'h40;
		memory[16'h2d57] <= 8'hdb;
		memory[16'h2d58] <= 8'hf5;
		memory[16'h2d59] <= 8'h6e;
		memory[16'h2d5a] <= 8'h79;
		memory[16'h2d5b] <= 8'hba;
		memory[16'h2d5c] <= 8'h74;
		memory[16'h2d5d] <= 8'h6b;
		memory[16'h2d5e] <= 8'h20;
		memory[16'h2d5f] <= 8'he3;
		memory[16'h2d60] <= 8'h40;
		memory[16'h2d61] <= 8'hb3;
		memory[16'h2d62] <= 8'h96;
		memory[16'h2d63] <= 8'h22;
		memory[16'h2d64] <= 8'h16;
		memory[16'h2d65] <= 8'hed;
		memory[16'h2d66] <= 8'h78;
		memory[16'h2d67] <= 8'h69;
		memory[16'h2d68] <= 8'hc5;
		memory[16'h2d69] <= 8'he5;
		memory[16'h2d6a] <= 8'h38;
		memory[16'h2d6b] <= 8'hce;
		memory[16'h2d6c] <= 8'h3c;
		memory[16'h2d6d] <= 8'h79;
		memory[16'h2d6e] <= 8'h1;
		memory[16'h2d6f] <= 8'hfa;
		memory[16'h2d70] <= 8'h30;
		memory[16'h2d71] <= 8'h11;
		memory[16'h2d72] <= 8'hb3;
		memory[16'h2d73] <= 8'h20;
		memory[16'h2d74] <= 8'h95;
		memory[16'h2d75] <= 8'hf3;
		memory[16'h2d76] <= 8'hfb;
		memory[16'h2d77] <= 8'h8a;
		memory[16'h2d78] <= 8'h61;
		memory[16'h2d79] <= 8'h74;
		memory[16'h2d7a] <= 8'h44;
		memory[16'h2d7b] <= 8'hd6;
		memory[16'h2d7c] <= 8'hdf;
		memory[16'h2d7d] <= 8'h64;
		memory[16'h2d7e] <= 8'hb9;
		memory[16'h2d7f] <= 8'h20;
		memory[16'h2d80] <= 8'h17;
		memory[16'h2d81] <= 8'h4f;
		memory[16'h2d82] <= 8'h42;
		memory[16'h2d83] <= 8'h2d;
		memory[16'h2d84] <= 8'h3d;
		memory[16'h2d85] <= 8'hba;
		memory[16'h2d86] <= 8'h97;
		memory[16'h2d87] <= 8'h2;
		memory[16'h2d88] <= 8'ha0;
		memory[16'h2d89] <= 8'hcf;
		memory[16'h2d8a] <= 8'hd1;
		memory[16'h2d8b] <= 8'hdc;
		memory[16'h2d8c] <= 8'h49;
		memory[16'h2d8d] <= 8'hd2;
		memory[16'h2d8e] <= 8'hd6;
		memory[16'h2d8f] <= 8'h79;
		memory[16'h2d90] <= 8'he3;
		memory[16'h2d91] <= 8'h89;
		memory[16'h2d92] <= 8'h99;
		memory[16'h2d93] <= 8'h78;
		memory[16'h2d94] <= 8'h7c;
		memory[16'h2d95] <= 8'h94;
		memory[16'h2d96] <= 8'h2;
		memory[16'h2d97] <= 8'hde;
		memory[16'h2d98] <= 8'h8;
		memory[16'h2d99] <= 8'h46;
		memory[16'h2d9a] <= 8'hb4;
		memory[16'h2d9b] <= 8'he8;
		memory[16'h2d9c] <= 8'haa;
		memory[16'h2d9d] <= 8'h6d;
		memory[16'h2d9e] <= 8'h8;
		memory[16'h2d9f] <= 8'hc1;
		memory[16'h2da0] <= 8'hbd;
		memory[16'h2da1] <= 8'h4a;
		memory[16'h2da2] <= 8'hee;
		memory[16'h2da3] <= 8'hfa;
		memory[16'h2da4] <= 8'h5;
		memory[16'h2da5] <= 8'h85;
		memory[16'h2da6] <= 8'hfc;
		memory[16'h2da7] <= 8'ha5;
		memory[16'h2da8] <= 8'h55;
		memory[16'h2da9] <= 8'hcd;
		memory[16'h2daa] <= 8'h81;
		memory[16'h2dab] <= 8'h9e;
		memory[16'h2dac] <= 8'h9f;
		memory[16'h2dad] <= 8'h58;
		memory[16'h2dae] <= 8'h17;
		memory[16'h2daf] <= 8'h82;
		memory[16'h2db0] <= 8'he1;
		memory[16'h2db1] <= 8'hb1;
		memory[16'h2db2] <= 8'hfa;
		memory[16'h2db3] <= 8'h5e;
		memory[16'h2db4] <= 8'h45;
		memory[16'h2db5] <= 8'hfc;
		memory[16'h2db6] <= 8'h3c;
		memory[16'h2db7] <= 8'h4e;
		memory[16'h2db8] <= 8'h42;
		memory[16'h2db9] <= 8'hf0;
		memory[16'h2dba] <= 8'h36;
		memory[16'h2dbb] <= 8'hec;
		memory[16'h2dbc] <= 8'h5d;
		memory[16'h2dbd] <= 8'h3e;
		memory[16'h2dbe] <= 8'had;
		memory[16'h2dbf] <= 8'h1a;
		memory[16'h2dc0] <= 8'h88;
		memory[16'h2dc1] <= 8'h9c;
		memory[16'h2dc2] <= 8'h14;
		memory[16'h2dc3] <= 8'h8d;
		memory[16'h2dc4] <= 8'h21;
		memory[16'h2dc5] <= 8'h11;
		memory[16'h2dc6] <= 8'h32;
		memory[16'h2dc7] <= 8'h76;
		memory[16'h2dc8] <= 8'hde;
		memory[16'h2dc9] <= 8'hb4;
		memory[16'h2dca] <= 8'h14;
		memory[16'h2dcb] <= 8'h7e;
		memory[16'h2dcc] <= 8'hc;
		memory[16'h2dcd] <= 8'h2c;
		memory[16'h2dce] <= 8'h0;
		memory[16'h2dcf] <= 8'hed;
		memory[16'h2dd0] <= 8'hdd;
		memory[16'h2dd1] <= 8'hfb;
		memory[16'h2dd2] <= 8'h4b;
		memory[16'h2dd3] <= 8'h22;
		memory[16'h2dd4] <= 8'hf7;
		memory[16'h2dd5] <= 8'h87;
		memory[16'h2dd6] <= 8'h70;
		memory[16'h2dd7] <= 8'h3a;
		memory[16'h2dd8] <= 8'h77;
		memory[16'h2dd9] <= 8'ha6;
		memory[16'h2dda] <= 8'h26;
		memory[16'h2ddb] <= 8'hd5;
		memory[16'h2ddc] <= 8'he4;
		memory[16'h2ddd] <= 8'hd4;
		memory[16'h2dde] <= 8'hef;
		memory[16'h2ddf] <= 8'h6d;
		memory[16'h2de0] <= 8'h70;
		memory[16'h2de1] <= 8'h4;
		memory[16'h2de2] <= 8'hfa;
		memory[16'h2de3] <= 8'h91;
		memory[16'h2de4] <= 8'h15;
		memory[16'h2de5] <= 8'h2d;
		memory[16'h2de6] <= 8'h8;
		memory[16'h2de7] <= 8'hf3;
		memory[16'h2de8] <= 8'he1;
		memory[16'h2de9] <= 8'h1c;
		memory[16'h2dea] <= 8'h71;
		memory[16'h2deb] <= 8'hed;
		memory[16'h2dec] <= 8'h48;
		memory[16'h2ded] <= 8'h72;
		memory[16'h2dee] <= 8'hda;
		memory[16'h2def] <= 8'h25;
		memory[16'h2df0] <= 8'h6d;
		memory[16'h2df1] <= 8'h26;
		memory[16'h2df2] <= 8'h48;
		memory[16'h2df3] <= 8'h64;
		memory[16'h2df4] <= 8'had;
		memory[16'h2df5] <= 8'hb8;
		memory[16'h2df6] <= 8'h9e;
		memory[16'h2df7] <= 8'h25;
		memory[16'h2df8] <= 8'h5f;
		memory[16'h2df9] <= 8'hc5;
		memory[16'h2dfa] <= 8'hfa;
		memory[16'h2dfb] <= 8'h43;
		memory[16'h2dfc] <= 8'h99;
		memory[16'h2dfd] <= 8'he9;
		memory[16'h2dfe] <= 8'hb0;
		memory[16'h2dff] <= 8'h9;
		memory[16'h2e00] <= 8'hed;
		memory[16'h2e01] <= 8'hab;
		memory[16'h2e02] <= 8'h9a;
		memory[16'h2e03] <= 8'h2;
		memory[16'h2e04] <= 8'hd8;
		memory[16'h2e05] <= 8'ha2;
		memory[16'h2e06] <= 8'hf6;
		memory[16'h2e07] <= 8'hb9;
		memory[16'h2e08] <= 8'hbf;
		memory[16'h2e09] <= 8'h67;
		memory[16'h2e0a] <= 8'ha6;
		memory[16'h2e0b] <= 8'h7;
		memory[16'h2e0c] <= 8'hd9;
		memory[16'h2e0d] <= 8'h80;
		memory[16'h2e0e] <= 8'h2d;
		memory[16'h2e0f] <= 8'h46;
		memory[16'h2e10] <= 8'ha6;
		memory[16'h2e11] <= 8'h75;
		memory[16'h2e12] <= 8'hab;
		memory[16'h2e13] <= 8'h54;
		memory[16'h2e14] <= 8'h2d;
		memory[16'h2e15] <= 8'h49;
		memory[16'h2e16] <= 8'h79;
		memory[16'h2e17] <= 8'h8c;
		memory[16'h2e18] <= 8'he;
		memory[16'h2e19] <= 8'h73;
		memory[16'h2e1a] <= 8'hd0;
		memory[16'h2e1b] <= 8'ha7;
		memory[16'h2e1c] <= 8'h5c;
		memory[16'h2e1d] <= 8'h80;
		memory[16'h2e1e] <= 8'hb0;
		memory[16'h2e1f] <= 8'h4a;
		memory[16'h2e20] <= 8'h2b;
		memory[16'h2e21] <= 8'h4b;
		memory[16'h2e22] <= 8'h4c;
		memory[16'h2e23] <= 8'h3;
		memory[16'h2e24] <= 8'hed;
		memory[16'h2e25] <= 8'h42;
		memory[16'h2e26] <= 8'hbc;
		memory[16'h2e27] <= 8'hac;
		memory[16'h2e28] <= 8'haa;
		memory[16'h2e29] <= 8'h62;
		memory[16'h2e2a] <= 8'hb4;
		memory[16'h2e2b] <= 8'h83;
		memory[16'h2e2c] <= 8'he3;
		memory[16'h2e2d] <= 8'he1;
		memory[16'h2e2e] <= 8'hca;
		memory[16'h2e2f] <= 8'h89;
		memory[16'h2e30] <= 8'h56;
		memory[16'h2e31] <= 8'h75;
		memory[16'h2e32] <= 8'hdd;
		memory[16'h2e33] <= 8'h83;
		memory[16'h2e34] <= 8'hbe;
		memory[16'h2e35] <= 8'h56;
		memory[16'h2e36] <= 8'h10;
		memory[16'h2e37] <= 8'hcd;
		memory[16'h2e38] <= 8'hc9;
		memory[16'h2e39] <= 8'he0;
		memory[16'h2e3a] <= 8'h74;
		memory[16'h2e3b] <= 8'h26;
		memory[16'h2e3c] <= 8'h60;
		memory[16'h2e3d] <= 8'h25;
		memory[16'h2e3e] <= 8'h70;
		memory[16'h2e3f] <= 8'h8c;
		memory[16'h2e40] <= 8'h70;
		memory[16'h2e41] <= 8'hbc;
		memory[16'h2e42] <= 8'h8f;
		memory[16'h2e43] <= 8'h5d;
		memory[16'h2e44] <= 8'hff;
		memory[16'h2e45] <= 8'h4c;
		memory[16'h2e46] <= 8'ha;
		memory[16'h2e47] <= 8'ha9;
		memory[16'h2e48] <= 8'hae;
		memory[16'h2e49] <= 8'hbe;
		memory[16'h2e4a] <= 8'h2c;
		memory[16'h2e4b] <= 8'h91;
		memory[16'h2e4c] <= 8'h9f;
		memory[16'h2e4d] <= 8'hf6;
		memory[16'h2e4e] <= 8'h1b;
		memory[16'h2e4f] <= 8'hf5;
		memory[16'h2e50] <= 8'h6b;
		memory[16'h2e51] <= 8'hf8;
		memory[16'h2e52] <= 8'h78;
		memory[16'h2e53] <= 8'h2a;
		memory[16'h2e54] <= 8'h4f;
		memory[16'h2e55] <= 8'h88;
		memory[16'h2e56] <= 8'hf7;
		memory[16'h2e57] <= 8'h18;
		memory[16'h2e58] <= 8'h68;
		memory[16'h2e59] <= 8'h6b;
		memory[16'h2e5a] <= 8'h3e;
		memory[16'h2e5b] <= 8'hc9;
		memory[16'h2e5c] <= 8'h90;
		memory[16'h2e5d] <= 8'hae;
		memory[16'h2e5e] <= 8'h55;
		memory[16'h2e5f] <= 8'h0;
		memory[16'h2e60] <= 8'h6b;
		memory[16'h2e61] <= 8'he4;
		memory[16'h2e62] <= 8'h5e;
		memory[16'h2e63] <= 8'h6a;
		memory[16'h2e64] <= 8'h30;
		memory[16'h2e65] <= 8'h68;
		memory[16'h2e66] <= 8'h13;
		memory[16'h2e67] <= 8'hdf;
		memory[16'h2e68] <= 8'h26;
		memory[16'h2e69] <= 8'h3f;
		memory[16'h2e6a] <= 8'h70;
		memory[16'h2e6b] <= 8'hc5;
		memory[16'h2e6c] <= 8'h36;
		memory[16'h2e6d] <= 8'h8b;
		memory[16'h2e6e] <= 8'hba;
		memory[16'h2e6f] <= 8'ha1;
		memory[16'h2e70] <= 8'h84;
		memory[16'h2e71] <= 8'h32;
		memory[16'h2e72] <= 8'hcb;
		memory[16'h2e73] <= 8'hd3;
		memory[16'h2e74] <= 8'hbb;
		memory[16'h2e75] <= 8'hc2;
		memory[16'h2e76] <= 8'heb;
		memory[16'h2e77] <= 8'h23;
		memory[16'h2e78] <= 8'h2e;
		memory[16'h2e79] <= 8'h2a;
		memory[16'h2e7a] <= 8'hec;
		memory[16'h2e7b] <= 8'hbe;
		memory[16'h2e7c] <= 8'hd8;
		memory[16'h2e7d] <= 8'h41;
		memory[16'h2e7e] <= 8'hbf;
		memory[16'h2e7f] <= 8'h43;
		memory[16'h2e80] <= 8'h26;
		memory[16'h2e81] <= 8'h1d;
		memory[16'h2e82] <= 8'had;
		memory[16'h2e83] <= 8'h56;
		memory[16'h2e84] <= 8'h85;
		memory[16'h2e85] <= 8'hc0;
		memory[16'h2e86] <= 8'h35;
		memory[16'h2e87] <= 8'hab;
		memory[16'h2e88] <= 8'h0;
		memory[16'h2e89] <= 8'ha6;
		memory[16'h2e8a] <= 8'h70;
		memory[16'h2e8b] <= 8'h36;
		memory[16'h2e8c] <= 8'h31;
		memory[16'h2e8d] <= 8'h2a;
		memory[16'h2e8e] <= 8'hd7;
		memory[16'h2e8f] <= 8'hb5;
		memory[16'h2e90] <= 8'h5c;
		memory[16'h2e91] <= 8'ha3;
		memory[16'h2e92] <= 8'h88;
		memory[16'h2e93] <= 8'h17;
		memory[16'h2e94] <= 8'h65;
		memory[16'h2e95] <= 8'h74;
		memory[16'h2e96] <= 8'h3b;
		memory[16'h2e97] <= 8'h93;
		memory[16'h2e98] <= 8'h9e;
		memory[16'h2e99] <= 8'h27;
		memory[16'h2e9a] <= 8'h52;
		memory[16'h2e9b] <= 8'h76;
		memory[16'h2e9c] <= 8'h69;
		memory[16'h2e9d] <= 8'h11;
		memory[16'h2e9e] <= 8'hba;
		memory[16'h2e9f] <= 8'h8f;
		memory[16'h2ea0] <= 8'h2e;
		memory[16'h2ea1] <= 8'h67;
		memory[16'h2ea2] <= 8'he5;
		memory[16'h2ea3] <= 8'hb3;
		memory[16'h2ea4] <= 8'h28;
		memory[16'h2ea5] <= 8'h1b;
		memory[16'h2ea6] <= 8'h5e;
		memory[16'h2ea7] <= 8'h28;
		memory[16'h2ea8] <= 8'hc1;
		memory[16'h2ea9] <= 8'hce;
		memory[16'h2eaa] <= 8'h5e;
		memory[16'h2eab] <= 8'hf2;
		memory[16'h2eac] <= 8'hf8;
		memory[16'h2ead] <= 8'h35;
		memory[16'h2eae] <= 8'ha8;
		memory[16'h2eaf] <= 8'h54;
		memory[16'h2eb0] <= 8'hd8;
		memory[16'h2eb1] <= 8'h30;
		memory[16'h2eb2] <= 8'h6c;
		memory[16'h2eb3] <= 8'h3e;
		memory[16'h2eb4] <= 8'ha4;
		memory[16'h2eb5] <= 8'ha7;
		memory[16'h2eb6] <= 8'hd1;
		memory[16'h2eb7] <= 8'h42;
		memory[16'h2eb8] <= 8'hce;
		memory[16'h2eb9] <= 8'h23;
		memory[16'h2eba] <= 8'hb9;
		memory[16'h2ebb] <= 8'h37;
		memory[16'h2ebc] <= 8'h34;
		memory[16'h2ebd] <= 8'h73;
		memory[16'h2ebe] <= 8'hc6;
		memory[16'h2ebf] <= 8'h62;
		memory[16'h2ec0] <= 8'hda;
		memory[16'h2ec1] <= 8'hac;
		memory[16'h2ec2] <= 8'h15;
		memory[16'h2ec3] <= 8'h2;
		memory[16'h2ec4] <= 8'hc7;
		memory[16'h2ec5] <= 8'h73;
		memory[16'h2ec6] <= 8'h2a;
		memory[16'h2ec7] <= 8'h88;
		memory[16'h2ec8] <= 8'h41;
		memory[16'h2ec9] <= 8'h88;
		memory[16'h2eca] <= 8'h7a;
		memory[16'h2ecb] <= 8'h39;
		memory[16'h2ecc] <= 8'hbe;
		memory[16'h2ecd] <= 8'h22;
		memory[16'h2ece] <= 8'h8e;
		memory[16'h2ecf] <= 8'h96;
		memory[16'h2ed0] <= 8'h53;
		memory[16'h2ed1] <= 8'hfa;
		memory[16'h2ed2] <= 8'hd4;
		memory[16'h2ed3] <= 8'hf7;
		memory[16'h2ed4] <= 8'ha1;
		memory[16'h2ed5] <= 8'ha6;
		memory[16'h2ed6] <= 8'h3a;
		memory[16'h2ed7] <= 8'h6f;
		memory[16'h2ed8] <= 8'hc9;
		memory[16'h2ed9] <= 8'hf3;
		memory[16'h2eda] <= 8'ha7;
		memory[16'h2edb] <= 8'hfe;
		memory[16'h2edc] <= 8'h66;
		memory[16'h2edd] <= 8'h6d;
		memory[16'h2ede] <= 8'h60;
		memory[16'h2edf] <= 8'h40;
		memory[16'h2ee0] <= 8'h19;
		memory[16'h2ee1] <= 8'h76;
		memory[16'h2ee2] <= 8'h43;
		memory[16'h2ee3] <= 8'he0;
		memory[16'h2ee4] <= 8'he9;
		memory[16'h2ee5] <= 8'h6d;
		memory[16'h2ee6] <= 8'h68;
		memory[16'h2ee7] <= 8'h2b;
		memory[16'h2ee8] <= 8'hf6;
		memory[16'h2ee9] <= 8'he3;
		memory[16'h2eea] <= 8'h64;
		memory[16'h2eeb] <= 8'hb4;
		memory[16'h2eec] <= 8'h5;
		memory[16'h2eed] <= 8'hf2;
		memory[16'h2eee] <= 8'h4a;
		memory[16'h2eef] <= 8'h58;
		memory[16'h2ef0] <= 8'hec;
		memory[16'h2ef1] <= 8'h1f;
		memory[16'h2ef2] <= 8'h50;
		memory[16'h2ef3] <= 8'h8d;
		memory[16'h2ef4] <= 8'hc5;
		memory[16'h2ef5] <= 8'h8a;
		memory[16'h2ef6] <= 8'hfd;
		memory[16'h2ef7] <= 8'h8e;
		memory[16'h2ef8] <= 8'h7d;
		memory[16'h2ef9] <= 8'ha4;
		memory[16'h2efa] <= 8'h8c;
		memory[16'h2efb] <= 8'he3;
		memory[16'h2efc] <= 8'h11;
		memory[16'h2efd] <= 8'hed;
		memory[16'h2efe] <= 8'h23;
		memory[16'h2eff] <= 8'h2b;
		memory[16'h2f00] <= 8'h63;
		memory[16'h2f01] <= 8'h66;
		memory[16'h2f02] <= 8'hb;
		memory[16'h2f03] <= 8'h4c;
		memory[16'h2f04] <= 8'hd4;
		memory[16'h2f05] <= 8'h74;
		memory[16'h2f06] <= 8'h77;
		memory[16'h2f07] <= 8'hca;
		memory[16'h2f08] <= 8'h57;
		memory[16'h2f09] <= 8'hdc;
		memory[16'h2f0a] <= 8'h7e;
		memory[16'h2f0b] <= 8'h5c;
		memory[16'h2f0c] <= 8'hce;
		memory[16'h2f0d] <= 8'hc8;
		memory[16'h2f0e] <= 8'hb5;
		memory[16'h2f0f] <= 8'hbb;
		memory[16'h2f10] <= 8'he7;
		memory[16'h2f11] <= 8'h5;
		memory[16'h2f12] <= 8'h48;
		memory[16'h2f13] <= 8'hac;
		memory[16'h2f14] <= 8'h8f;
		memory[16'h2f15] <= 8'h45;
		memory[16'h2f16] <= 8'h3b;
		memory[16'h2f17] <= 8'hc;
		memory[16'h2f18] <= 8'he9;
		memory[16'h2f19] <= 8'hc7;
		memory[16'h2f1a] <= 8'hef;
		memory[16'h2f1b] <= 8'hfb;
		memory[16'h2f1c] <= 8'hb4;
		memory[16'h2f1d] <= 8'h12;
		memory[16'h2f1e] <= 8'h26;
		memory[16'h2f1f] <= 8'h17;
		memory[16'h2f20] <= 8'h79;
		memory[16'h2f21] <= 8'h31;
		memory[16'h2f22] <= 8'h64;
		memory[16'h2f23] <= 8'h4d;
		memory[16'h2f24] <= 8'ha5;
		memory[16'h2f25] <= 8'hdb;
		memory[16'h2f26] <= 8'h17;
		memory[16'h2f27] <= 8'hfc;
		memory[16'h2f28] <= 8'hb7;
		memory[16'h2f29] <= 8'h95;
		memory[16'h2f2a] <= 8'h59;
		memory[16'h2f2b] <= 8'h86;
		memory[16'h2f2c] <= 8'h5d;
		memory[16'h2f2d] <= 8'he;
		memory[16'h2f2e] <= 8'h41;
		memory[16'h2f2f] <= 8'h45;
		memory[16'h2f30] <= 8'h13;
		memory[16'h2f31] <= 8'h89;
		memory[16'h2f32] <= 8'hf1;
		memory[16'h2f33] <= 8'ha2;
		memory[16'h2f34] <= 8'hcf;
		memory[16'h2f35] <= 8'h2c;
		memory[16'h2f36] <= 8'hae;
		memory[16'h2f37] <= 8'hb8;
		memory[16'h2f38] <= 8'hf4;
		memory[16'h2f39] <= 8'h9d;
		memory[16'h2f3a] <= 8'hb3;
		memory[16'h2f3b] <= 8'ha8;
		memory[16'h2f3c] <= 8'haf;
		memory[16'h2f3d] <= 8'hd9;
		memory[16'h2f3e] <= 8'hc0;
		memory[16'h2f3f] <= 8'h28;
		memory[16'h2f40] <= 8'hb;
		memory[16'h2f41] <= 8'h24;
		memory[16'h2f42] <= 8'h75;
		memory[16'h2f43] <= 8'hb0;
		memory[16'h2f44] <= 8'hff;
		memory[16'h2f45] <= 8'h8c;
		memory[16'h2f46] <= 8'had;
		memory[16'h2f47] <= 8'hb7;
		memory[16'h2f48] <= 8'h21;
		memory[16'h2f49] <= 8'h6;
		memory[16'h2f4a] <= 8'h3d;
		memory[16'h2f4b] <= 8'h7f;
		memory[16'h2f4c] <= 8'h14;
		memory[16'h2f4d] <= 8'h7e;
		memory[16'h2f4e] <= 8'hc4;
		memory[16'h2f4f] <= 8'h27;
		memory[16'h2f50] <= 8'h7;
		memory[16'h2f51] <= 8'hb5;
		memory[16'h2f52] <= 8'hc9;
		memory[16'h2f53] <= 8'hd6;
		memory[16'h2f54] <= 8'he2;
		memory[16'h2f55] <= 8'h77;
		memory[16'h2f56] <= 8'h8f;
		memory[16'h2f57] <= 8'hd6;
		memory[16'h2f58] <= 8'h14;
		memory[16'h2f59] <= 8'h42;
		memory[16'h2f5a] <= 8'h7e;
		memory[16'h2f5b] <= 8'hc3;
		memory[16'h2f5c] <= 8'h1c;
		memory[16'h2f5d] <= 8'h3e;
		memory[16'h2f5e] <= 8'hec;
		memory[16'h2f5f] <= 8'h27;
		memory[16'h2f60] <= 8'h62;
		memory[16'h2f61] <= 8'h61;
		memory[16'h2f62] <= 8'hd7;
		memory[16'h2f63] <= 8'h62;
		memory[16'h2f64] <= 8'hee;
		memory[16'h2f65] <= 8'h84;
		memory[16'h2f66] <= 8'h19;
		memory[16'h2f67] <= 8'hf;
		memory[16'h2f68] <= 8'h8a;
		memory[16'h2f69] <= 8'h56;
		memory[16'h2f6a] <= 8'h8e;
		memory[16'h2f6b] <= 8'h9e;
		memory[16'h2f6c] <= 8'hd4;
		memory[16'h2f6d] <= 8'h52;
		memory[16'h2f6e] <= 8'hc5;
		memory[16'h2f6f] <= 8'hdb;
		memory[16'h2f70] <= 8'h8;
		memory[16'h2f71] <= 8'h8e;
		memory[16'h2f72] <= 8'hb2;
		memory[16'h2f73] <= 8'hea;
		memory[16'h2f74] <= 8'h5;
		memory[16'h2f75] <= 8'h41;
		memory[16'h2f76] <= 8'hc0;
		memory[16'h2f77] <= 8'h19;
		memory[16'h2f78] <= 8'h83;
		memory[16'h2f79] <= 8'h3e;
		memory[16'h2f7a] <= 8'hdd;
		memory[16'h2f7b] <= 8'h9f;
		memory[16'h2f7c] <= 8'h7d;
		memory[16'h2f7d] <= 8'hc9;
		memory[16'h2f7e] <= 8'hc6;
		memory[16'h2f7f] <= 8'hdf;
		memory[16'h2f80] <= 8'h2a;
		memory[16'h2f81] <= 8'h9e;
		memory[16'h2f82] <= 8'h41;
		memory[16'h2f83] <= 8'h18;
		memory[16'h2f84] <= 8'h22;
		memory[16'h2f85] <= 8'h5a;
		memory[16'h2f86] <= 8'h28;
		memory[16'h2f87] <= 8'had;
		memory[16'h2f88] <= 8'hb0;
		memory[16'h2f89] <= 8'hb6;
		memory[16'h2f8a] <= 8'h4b;
		memory[16'h2f8b] <= 8'h84;
		memory[16'h2f8c] <= 8'h9;
		memory[16'h2f8d] <= 8'h11;
		memory[16'h2f8e] <= 8'h60;
		memory[16'h2f8f] <= 8'h11;
		memory[16'h2f90] <= 8'h9f;
		memory[16'h2f91] <= 8'h12;
		memory[16'h2f92] <= 8'hfb;
		memory[16'h2f93] <= 8'ha5;
		memory[16'h2f94] <= 8'h53;
		memory[16'h2f95] <= 8'hbb;
		memory[16'h2f96] <= 8'hbe;
		memory[16'h2f97] <= 8'hd6;
		memory[16'h2f98] <= 8'hf9;
		memory[16'h2f99] <= 8'h9b;
		memory[16'h2f9a] <= 8'h76;
		memory[16'h2f9b] <= 8'h76;
		memory[16'h2f9c] <= 8'h64;
		memory[16'h2f9d] <= 8'h3c;
		memory[16'h2f9e] <= 8'h56;
		memory[16'h2f9f] <= 8'h8f;
		memory[16'h2fa0] <= 8'hda;
		memory[16'h2fa1] <= 8'h97;
		memory[16'h2fa2] <= 8'ha7;
		memory[16'h2fa3] <= 8'hfd;
		memory[16'h2fa4] <= 8'hf2;
		memory[16'h2fa5] <= 8'hcf;
		memory[16'h2fa6] <= 8'haa;
		memory[16'h2fa7] <= 8'ha2;
		memory[16'h2fa8] <= 8'h86;
		memory[16'h2fa9] <= 8'hf5;
		memory[16'h2faa] <= 8'h27;
		memory[16'h2fab] <= 8'h8f;
		memory[16'h2fac] <= 8'h6;
		memory[16'h2fad] <= 8'h87;
		memory[16'h2fae] <= 8'ha0;
		memory[16'h2faf] <= 8'ha6;
		memory[16'h2fb0] <= 8'h99;
		memory[16'h2fb1] <= 8'h9b;
		memory[16'h2fb2] <= 8'h4b;
		memory[16'h2fb3] <= 8'hec;
		memory[16'h2fb4] <= 8'h56;
		memory[16'h2fb5] <= 8'h9;
		memory[16'h2fb6] <= 8'hc2;
		memory[16'h2fb7] <= 8'h4f;
		memory[16'h2fb8] <= 8'ha5;
		memory[16'h2fb9] <= 8'h38;
		memory[16'h2fba] <= 8'hc6;
		memory[16'h2fbb] <= 8'h9;
		memory[16'h2fbc] <= 8'h75;
		memory[16'h2fbd] <= 8'h1c;
		memory[16'h2fbe] <= 8'h98;
		memory[16'h2fbf] <= 8'h4f;
		memory[16'h2fc0] <= 8'hb3;
		memory[16'h2fc1] <= 8'h40;
		memory[16'h2fc2] <= 8'h4c;
		memory[16'h2fc3] <= 8'ha5;
		memory[16'h2fc4] <= 8'hf;
		memory[16'h2fc5] <= 8'hf6;
		memory[16'h2fc6] <= 8'h48;
		memory[16'h2fc7] <= 8'h95;
		memory[16'h2fc8] <= 8'hec;
		memory[16'h2fc9] <= 8'h6f;
		memory[16'h2fca] <= 8'h24;
		memory[16'h2fcb] <= 8'hf2;
		memory[16'h2fcc] <= 8'hf6;
		memory[16'h2fcd] <= 8'hc4;
		memory[16'h2fce] <= 8'h98;
		memory[16'h2fcf] <= 8'h8f;
		memory[16'h2fd0] <= 8'h5f;
		memory[16'h2fd1] <= 8'he3;
		memory[16'h2fd2] <= 8'h7b;
		memory[16'h2fd3] <= 8'hb5;
		memory[16'h2fd4] <= 8'hed;
		memory[16'h2fd5] <= 8'h3d;
		memory[16'h2fd6] <= 8'h5;
		memory[16'h2fd7] <= 8'h92;
		memory[16'h2fd8] <= 8'h76;
		memory[16'h2fd9] <= 8'hcb;
		memory[16'h2fda] <= 8'h9b;
		memory[16'h2fdb] <= 8'heb;
		memory[16'h2fdc] <= 8'he7;
		memory[16'h2fdd] <= 8'h34;
		memory[16'h2fde] <= 8'h3a;
		memory[16'h2fdf] <= 8'h9a;
		memory[16'h2fe0] <= 8'h74;
		memory[16'h2fe1] <= 8'h87;
		memory[16'h2fe2] <= 8'h40;
		memory[16'h2fe3] <= 8'h83;
		memory[16'h2fe4] <= 8'h7d;
		memory[16'h2fe5] <= 8'h88;
		memory[16'h2fe6] <= 8'h19;
		memory[16'h2fe7] <= 8'h69;
		memory[16'h2fe8] <= 8'hf7;
		memory[16'h2fe9] <= 8'h3d;
		memory[16'h2fea] <= 8'h5c;
		memory[16'h2feb] <= 8'hed;
		memory[16'h2fec] <= 8'h2;
		memory[16'h2fed] <= 8'hf4;
		memory[16'h2fee] <= 8'h7c;
		memory[16'h2fef] <= 8'h61;
		memory[16'h2ff0] <= 8'hd8;
		memory[16'h2ff1] <= 8'hf7;
		memory[16'h2ff2] <= 8'h17;
		memory[16'h2ff3] <= 8'hc5;
		memory[16'h2ff4] <= 8'h34;
		memory[16'h2ff5] <= 8'h1c;
		memory[16'h2ff6] <= 8'h57;
		memory[16'h2ff7] <= 8'haa;
		memory[16'h2ff8] <= 8'he7;
		memory[16'h2ff9] <= 8'hf2;
		memory[16'h2ffa] <= 8'h95;
		memory[16'h2ffb] <= 8'hce;
		memory[16'h2ffc] <= 8'h26;
		memory[16'h2ffd] <= 8'hd0;
		memory[16'h2ffe] <= 8'h68;
		memory[16'h2fff] <= 8'h9a;
		memory[16'h3000] <= 8'h57;
		memory[16'h3001] <= 8'ha8;
		memory[16'h3002] <= 8'h1e;
		memory[16'h3003] <= 8'hd4;
		memory[16'h3004] <= 8'h30;
		memory[16'h3005] <= 8'h37;
		memory[16'h3006] <= 8'h3e;
		memory[16'h3007] <= 8'h27;
		memory[16'h3008] <= 8'h74;
		memory[16'h3009] <= 8'h9a;
		memory[16'h300a] <= 8'h14;
		memory[16'h300b] <= 8'h76;
		memory[16'h300c] <= 8'h8e;
		memory[16'h300d] <= 8'h90;
		memory[16'h300e] <= 8'hd8;
		memory[16'h300f] <= 8'h66;
		memory[16'h3010] <= 8'h87;
		memory[16'h3011] <= 8'hef;
		memory[16'h3012] <= 8'h2b;
		memory[16'h3013] <= 8'hbc;
		memory[16'h3014] <= 8'hb;
		memory[16'h3015] <= 8'h82;
		memory[16'h3016] <= 8'h66;
		memory[16'h3017] <= 8'hf2;
		memory[16'h3018] <= 8'h75;
		memory[16'h3019] <= 8'hfc;
		memory[16'h301a] <= 8'hc0;
		memory[16'h301b] <= 8'h9b;
		memory[16'h301c] <= 8'hcc;
		memory[16'h301d] <= 8'h28;
		memory[16'h301e] <= 8'h36;
		memory[16'h301f] <= 8'h23;
		memory[16'h3020] <= 8'hd1;
		memory[16'h3021] <= 8'h54;
		memory[16'h3022] <= 8'hf7;
		memory[16'h3023] <= 8'h1;
		memory[16'h3024] <= 8'h8b;
		memory[16'h3025] <= 8'h35;
		memory[16'h3026] <= 8'h29;
		memory[16'h3027] <= 8'hff;
		memory[16'h3028] <= 8'hcf;
		memory[16'h3029] <= 8'h3d;
		memory[16'h302a] <= 8'h76;
		memory[16'h302b] <= 8'h5e;
		memory[16'h302c] <= 8'hce;
		memory[16'h302d] <= 8'h4e;
		memory[16'h302e] <= 8'hc4;
		memory[16'h302f] <= 8'h55;
		memory[16'h3030] <= 8'h3d;
		memory[16'h3031] <= 8'hf0;
		memory[16'h3032] <= 8'h11;
		memory[16'h3033] <= 8'h48;
		memory[16'h3034] <= 8'h72;
		memory[16'h3035] <= 8'h78;
		memory[16'h3036] <= 8'h3a;
		memory[16'h3037] <= 8'he7;
		memory[16'h3038] <= 8'h74;
		memory[16'h3039] <= 8'hfa;
		memory[16'h303a] <= 8'h83;
		memory[16'h303b] <= 8'h40;
		memory[16'h303c] <= 8'h22;
		memory[16'h303d] <= 8'hb9;
		memory[16'h303e] <= 8'h63;
		memory[16'h303f] <= 8'hf3;
		memory[16'h3040] <= 8'hd;
		memory[16'h3041] <= 8'h5a;
		memory[16'h3042] <= 8'hf5;
		memory[16'h3043] <= 8'h98;
		memory[16'h3044] <= 8'h90;
		memory[16'h3045] <= 8'h1e;
		memory[16'h3046] <= 8'h97;
		memory[16'h3047] <= 8'h5f;
		memory[16'h3048] <= 8'h5b;
		memory[16'h3049] <= 8'hd;
		memory[16'h304a] <= 8'hbd;
		memory[16'h304b] <= 8'h29;
		memory[16'h304c] <= 8'h5b;
		memory[16'h304d] <= 8'h82;
		memory[16'h304e] <= 8'h7f;
		memory[16'h304f] <= 8'h98;
		memory[16'h3050] <= 8'h72;
		memory[16'h3051] <= 8'h90;
		memory[16'h3052] <= 8'he0;
		memory[16'h3053] <= 8'he4;
		memory[16'h3054] <= 8'h8;
		memory[16'h3055] <= 8'h1a;
		memory[16'h3056] <= 8'hcc;
		memory[16'h3057] <= 8'h7c;
		memory[16'h3058] <= 8'h14;
		memory[16'h3059] <= 8'h4f;
		memory[16'h305a] <= 8'hbc;
		memory[16'h305b] <= 8'h37;
		memory[16'h305c] <= 8'h8;
		memory[16'h305d] <= 8'h1f;
		memory[16'h305e] <= 8'h2a;
		memory[16'h305f] <= 8'h15;
		memory[16'h3060] <= 8'h7a;
		memory[16'h3061] <= 8'h1f;
		memory[16'h3062] <= 8'had;
		memory[16'h3063] <= 8'ha;
		memory[16'h3064] <= 8'h3d;
		memory[16'h3065] <= 8'h44;
		memory[16'h3066] <= 8'h69;
		memory[16'h3067] <= 8'h99;
		memory[16'h3068] <= 8'h52;
		memory[16'h3069] <= 8'h27;
		memory[16'h306a] <= 8'hc2;
		memory[16'h306b] <= 8'had;
		memory[16'h306c] <= 8'ha9;
		memory[16'h306d] <= 8'h41;
		memory[16'h306e] <= 8'h46;
		memory[16'h306f] <= 8'h1b;
		memory[16'h3070] <= 8'hd2;
		memory[16'h3071] <= 8'h26;
		memory[16'h3072] <= 8'hff;
		memory[16'h3073] <= 8'hda;
		memory[16'h3074] <= 8'h41;
		memory[16'h3075] <= 8'hcb;
		memory[16'h3076] <= 8'h57;
		memory[16'h3077] <= 8'h55;
		memory[16'h3078] <= 8'h1a;
		memory[16'h3079] <= 8'h13;
		memory[16'h307a] <= 8'h8c;
		memory[16'h307b] <= 8'h22;
		memory[16'h307c] <= 8'h33;
		memory[16'h307d] <= 8'hb7;
		memory[16'h307e] <= 8'h37;
		memory[16'h307f] <= 8'had;
		memory[16'h3080] <= 8'hd6;
		memory[16'h3081] <= 8'he4;
		memory[16'h3082] <= 8'hb7;
		memory[16'h3083] <= 8'h14;
		memory[16'h3084] <= 8'h29;
		memory[16'h3085] <= 8'h20;
		memory[16'h3086] <= 8'had;
		memory[16'h3087] <= 8'h7b;
		memory[16'h3088] <= 8'h47;
		memory[16'h3089] <= 8'h6f;
		memory[16'h308a] <= 8'h28;
		memory[16'h308b] <= 8'hf0;
		memory[16'h308c] <= 8'hb1;
		memory[16'h308d] <= 8'h6e;
		memory[16'h308e] <= 8'hb;
		memory[16'h308f] <= 8'h83;
		memory[16'h3090] <= 8'h95;
		memory[16'h3091] <= 8'hb;
		memory[16'h3092] <= 8'h5d;
		memory[16'h3093] <= 8'hd6;
		memory[16'h3094] <= 8'hd6;
		memory[16'h3095] <= 8'hb4;
		memory[16'h3096] <= 8'h2b;
		memory[16'h3097] <= 8'hf1;
		memory[16'h3098] <= 8'hc8;
		memory[16'h3099] <= 8'hb8;
		memory[16'h309a] <= 8'h13;
		memory[16'h309b] <= 8'hfb;
		memory[16'h309c] <= 8'h6f;
		memory[16'h309d] <= 8'h4b;
		memory[16'h309e] <= 8'ha8;
		memory[16'h309f] <= 8'h45;
		memory[16'h30a0] <= 8'h2f;
		memory[16'h30a1] <= 8'h5f;
		memory[16'h30a2] <= 8'h59;
		memory[16'h30a3] <= 8'h58;
		memory[16'h30a4] <= 8'h7f;
		memory[16'h30a5] <= 8'h6;
		memory[16'h30a6] <= 8'hd3;
		memory[16'h30a7] <= 8'hc7;
		memory[16'h30a8] <= 8'h76;
		memory[16'h30a9] <= 8'hfc;
		memory[16'h30aa] <= 8'hb7;
		memory[16'h30ab] <= 8'h27;
		memory[16'h30ac] <= 8'h6a;
		memory[16'h30ad] <= 8'hc3;
		memory[16'h30ae] <= 8'haa;
		memory[16'h30af] <= 8'hff;
		memory[16'h30b0] <= 8'hce;
		memory[16'h30b1] <= 8'h7;
		memory[16'h30b2] <= 8'hd5;
		memory[16'h30b3] <= 8'ha4;
		memory[16'h30b4] <= 8'hbc;
		memory[16'h30b5] <= 8'h1;
		memory[16'h30b6] <= 8'h95;
		memory[16'h30b7] <= 8'h84;
		memory[16'h30b8] <= 8'hb9;
		memory[16'h30b9] <= 8'ha9;
		memory[16'h30ba] <= 8'h7f;
		memory[16'h30bb] <= 8'h28;
		memory[16'h30bc] <= 8'hf4;
		memory[16'h30bd] <= 8'h27;
		memory[16'h30be] <= 8'h6d;
		memory[16'h30bf] <= 8'h23;
		memory[16'h30c0] <= 8'h86;
		memory[16'h30c1] <= 8'hc7;
		memory[16'h30c2] <= 8'h7c;
		memory[16'h30c3] <= 8'h5;
		memory[16'h30c4] <= 8'hcd;
		memory[16'h30c5] <= 8'h4f;
		memory[16'h30c6] <= 8'hcc;
		memory[16'h30c7] <= 8'h43;
		memory[16'h30c8] <= 8'h4b;
		memory[16'h30c9] <= 8'h84;
		memory[16'h30ca] <= 8'h6a;
		memory[16'h30cb] <= 8'hb6;
		memory[16'h30cc] <= 8'h47;
		memory[16'h30cd] <= 8'h14;
		memory[16'h30ce] <= 8'hb5;
		memory[16'h30cf] <= 8'h15;
		memory[16'h30d0] <= 8'h1c;
		memory[16'h30d1] <= 8'h8b;
		memory[16'h30d2] <= 8'hb9;
		memory[16'h30d3] <= 8'hd8;
		memory[16'h30d4] <= 8'h8c;
		memory[16'h30d5] <= 8'h4f;
		memory[16'h30d6] <= 8'h5c;
		memory[16'h30d7] <= 8'h45;
		memory[16'h30d8] <= 8'hf8;
		memory[16'h30d9] <= 8'hdb;
		memory[16'h30da] <= 8'h6d;
		memory[16'h30db] <= 8'hec;
		memory[16'h30dc] <= 8'h2;
		memory[16'h30dd] <= 8'hda;
		memory[16'h30de] <= 8'hf;
		memory[16'h30df] <= 8'h88;
		memory[16'h30e0] <= 8'ha1;
		memory[16'h30e1] <= 8'h8b;
		memory[16'h30e2] <= 8'h8d;
		memory[16'h30e3] <= 8'h6f;
		memory[16'h30e4] <= 8'hdb;
		memory[16'h30e5] <= 8'h5a;
		memory[16'h30e6] <= 8'hb2;
		memory[16'h30e7] <= 8'h26;
		memory[16'h30e8] <= 8'hde;
		memory[16'h30e9] <= 8'h1d;
		memory[16'h30ea] <= 8'hdc;
		memory[16'h30eb] <= 8'h25;
		memory[16'h30ec] <= 8'h31;
		memory[16'h30ed] <= 8'h92;
		memory[16'h30ee] <= 8'h3a;
		memory[16'h30ef] <= 8'h4d;
		memory[16'h30f0] <= 8'h1d;
		memory[16'h30f1] <= 8'hf3;
		memory[16'h30f2] <= 8'h25;
		memory[16'h30f3] <= 8'ha9;
		memory[16'h30f4] <= 8'h42;
		memory[16'h30f5] <= 8'h81;
		memory[16'h30f6] <= 8'hee;
		memory[16'h30f7] <= 8'h3a;
		memory[16'h30f8] <= 8'h5c;
		memory[16'h30f9] <= 8'h5b;
		memory[16'h30fa] <= 8'h26;
		memory[16'h30fb] <= 8'h5e;
		memory[16'h30fc] <= 8'h35;
		memory[16'h30fd] <= 8'h36;
		memory[16'h30fe] <= 8'he6;
		memory[16'h30ff] <= 8'hd7;
		memory[16'h3100] <= 8'hc1;
		memory[16'h3101] <= 8'h74;
		memory[16'h3102] <= 8'h46;
		memory[16'h3103] <= 8'h9c;
		memory[16'h3104] <= 8'hce;
		memory[16'h3105] <= 8'hf8;
		memory[16'h3106] <= 8'hc3;
		memory[16'h3107] <= 8'hac;
		memory[16'h3108] <= 8'h15;
		memory[16'h3109] <= 8'h9f;
		memory[16'h310a] <= 8'hd1;
		memory[16'h310b] <= 8'h47;
		memory[16'h310c] <= 8'h31;
		memory[16'h310d] <= 8'hb;
		memory[16'h310e] <= 8'h94;
		memory[16'h310f] <= 8'h4e;
		memory[16'h3110] <= 8'hfe;
		memory[16'h3111] <= 8'hba;
		memory[16'h3112] <= 8'hf7;
		memory[16'h3113] <= 8'h41;
		memory[16'h3114] <= 8'h3b;
		memory[16'h3115] <= 8'he5;
		memory[16'h3116] <= 8'h7b;
		memory[16'h3117] <= 8'h98;
		memory[16'h3118] <= 8'h40;
		memory[16'h3119] <= 8'ha2;
		memory[16'h311a] <= 8'hf6;
		memory[16'h311b] <= 8'h76;
		memory[16'h311c] <= 8'hd8;
		memory[16'h311d] <= 8'hdd;
		memory[16'h311e] <= 8'h4d;
		memory[16'h311f] <= 8'h99;
		memory[16'h3120] <= 8'h51;
		memory[16'h3121] <= 8'h93;
		memory[16'h3122] <= 8'h36;
		memory[16'h3123] <= 8'h1f;
		memory[16'h3124] <= 8'h8b;
		memory[16'h3125] <= 8'hf9;
		memory[16'h3126] <= 8'hcb;
		memory[16'h3127] <= 8'ha1;
		memory[16'h3128] <= 8'h98;
		memory[16'h3129] <= 8'h9c;
		memory[16'h312a] <= 8'he8;
		memory[16'h312b] <= 8'hca;
		memory[16'h312c] <= 8'ha7;
		memory[16'h312d] <= 8'h7c;
		memory[16'h312e] <= 8'h18;
		memory[16'h312f] <= 8'ha5;
		memory[16'h3130] <= 8'h36;
		memory[16'h3131] <= 8'h10;
		memory[16'h3132] <= 8'he6;
		memory[16'h3133] <= 8'h72;
		memory[16'h3134] <= 8'hf5;
		memory[16'h3135] <= 8'h62;
		memory[16'h3136] <= 8'ha;
		memory[16'h3137] <= 8'h36;
		memory[16'h3138] <= 8'h4;
		memory[16'h3139] <= 8'h0;
		memory[16'h313a] <= 8'hac;
		memory[16'h313b] <= 8'hdc;
		memory[16'h313c] <= 8'hdd;
		memory[16'h313d] <= 8'hf9;
		memory[16'h313e] <= 8'h75;
		memory[16'h313f] <= 8'h2e;
		memory[16'h3140] <= 8'h8c;
		memory[16'h3141] <= 8'hab;
		memory[16'h3142] <= 8'h4d;
		memory[16'h3143] <= 8'h17;
		memory[16'h3144] <= 8'ha4;
		memory[16'h3145] <= 8'h18;
		memory[16'h3146] <= 8'hb8;
		memory[16'h3147] <= 8'h3d;
		memory[16'h3148] <= 8'hb4;
		memory[16'h3149] <= 8'ha0;
		memory[16'h314a] <= 8'h7;
		memory[16'h314b] <= 8'h5b;
		memory[16'h314c] <= 8'h1d;
		memory[16'h314d] <= 8'h1f;
		memory[16'h314e] <= 8'h1;
		memory[16'h314f] <= 8'h53;
		memory[16'h3150] <= 8'h2f;
		memory[16'h3151] <= 8'he7;
		memory[16'h3152] <= 8'hc5;
		memory[16'h3153] <= 8'h25;
		memory[16'h3154] <= 8'h49;
		memory[16'h3155] <= 8'hcf;
		memory[16'h3156] <= 8'h5b;
		memory[16'h3157] <= 8'h4d;
		memory[16'h3158] <= 8'hd0;
		memory[16'h3159] <= 8'h7;
		memory[16'h315a] <= 8'h29;
		memory[16'h315b] <= 8'had;
		memory[16'h315c] <= 8'h0;
		memory[16'h315d] <= 8'h9f;
		memory[16'h315e] <= 8'hdc;
		memory[16'h315f] <= 8'h8c;
		memory[16'h3160] <= 8'h4a;
		memory[16'h3161] <= 8'h29;
		memory[16'h3162] <= 8'ha3;
		memory[16'h3163] <= 8'hef;
		memory[16'h3164] <= 8'h42;
		memory[16'h3165] <= 8'h5c;
		memory[16'h3166] <= 8'h2c;
		memory[16'h3167] <= 8'hf6;
		memory[16'h3168] <= 8'hfc;
		memory[16'h3169] <= 8'h33;
		memory[16'h316a] <= 8'h52;
		memory[16'h316b] <= 8'h19;
		memory[16'h316c] <= 8'h52;
		memory[16'h316d] <= 8'h53;
		memory[16'h316e] <= 8'h6d;
		memory[16'h316f] <= 8'h82;
		memory[16'h3170] <= 8'h3a;
		memory[16'h3171] <= 8'h32;
		memory[16'h3172] <= 8'ha7;
		memory[16'h3173] <= 8'h84;
		memory[16'h3174] <= 8'h2;
		memory[16'h3175] <= 8'h2;
		memory[16'h3176] <= 8'hd1;
		memory[16'h3177] <= 8'hd2;
		memory[16'h3178] <= 8'h9;
		memory[16'h3179] <= 8'hfb;
		memory[16'h317a] <= 8'h7f;
		memory[16'h317b] <= 8'h9;
		memory[16'h317c] <= 8'h9a;
		memory[16'h317d] <= 8'h5b;
		memory[16'h317e] <= 8'h95;
		memory[16'h317f] <= 8'he4;
		memory[16'h3180] <= 8'h85;
		memory[16'h3181] <= 8'h38;
		memory[16'h3182] <= 8'hd3;
		memory[16'h3183] <= 8'hc7;
		memory[16'h3184] <= 8'h94;
		memory[16'h3185] <= 8'hff;
		memory[16'h3186] <= 8'hbd;
		memory[16'h3187] <= 8'h91;
		memory[16'h3188] <= 8'h32;
		memory[16'h3189] <= 8'hf;
		memory[16'h318a] <= 8'haa;
		memory[16'h318b] <= 8'h85;
		memory[16'h318c] <= 8'h62;
		memory[16'h318d] <= 8'h17;
		memory[16'h318e] <= 8'h7;
		memory[16'h318f] <= 8'h9d;
		memory[16'h3190] <= 8'h4a;
		memory[16'h3191] <= 8'hae;
		memory[16'h3192] <= 8'h21;
		memory[16'h3193] <= 8'h4c;
		memory[16'h3194] <= 8'hb0;
		memory[16'h3195] <= 8'hf2;
		memory[16'h3196] <= 8'h1e;
		memory[16'h3197] <= 8'hb9;
		memory[16'h3198] <= 8'hed;
		memory[16'h3199] <= 8'h9d;
		memory[16'h319a] <= 8'hc2;
		memory[16'h319b] <= 8'h87;
		memory[16'h319c] <= 8'hf9;
		memory[16'h319d] <= 8'h57;
		memory[16'h319e] <= 8'h6c;
		memory[16'h319f] <= 8'h7e;
		memory[16'h31a0] <= 8'h8f;
		memory[16'h31a1] <= 8'h3f;
		memory[16'h31a2] <= 8'h45;
		memory[16'h31a3] <= 8'h24;
		memory[16'h31a4] <= 8'h3f;
		memory[16'h31a5] <= 8'h2;
		memory[16'h31a6] <= 8'hb5;
		memory[16'h31a7] <= 8'h71;
		memory[16'h31a8] <= 8'h12;
		memory[16'h31a9] <= 8'h5f;
		memory[16'h31aa] <= 8'hf6;
		memory[16'h31ab] <= 8'h74;
		memory[16'h31ac] <= 8'h77;
		memory[16'h31ad] <= 8'hfd;
		memory[16'h31ae] <= 8'h11;
		memory[16'h31af] <= 8'hc1;
		memory[16'h31b0] <= 8'hab;
		memory[16'h31b1] <= 8'h32;
		memory[16'h31b2] <= 8'hd;
		memory[16'h31b3] <= 8'h5b;
		memory[16'h31b4] <= 8'h25;
		memory[16'h31b5] <= 8'h2b;
		memory[16'h31b6] <= 8'h14;
		memory[16'h31b7] <= 8'h12;
		memory[16'h31b8] <= 8'hc8;
		memory[16'h31b9] <= 8'hd6;
		memory[16'h31ba] <= 8'h9a;
		memory[16'h31bb] <= 8'hc1;
		memory[16'h31bc] <= 8'h2d;
		memory[16'h31bd] <= 8'h6;
		memory[16'h31be] <= 8'h3f;
		memory[16'h31bf] <= 8'hbd;
		memory[16'h31c0] <= 8'h45;
		memory[16'h31c1] <= 8'h84;
		memory[16'h31c2] <= 8'he1;
		memory[16'h31c3] <= 8'h84;
		memory[16'h31c4] <= 8'h87;
		memory[16'h31c5] <= 8'h96;
		memory[16'h31c6] <= 8'hf6;
		memory[16'h31c7] <= 8'h99;
		memory[16'h31c8] <= 8'hf5;
		memory[16'h31c9] <= 8'hec;
		memory[16'h31ca] <= 8'hd;
		memory[16'h31cb] <= 8'h6c;
		memory[16'h31cc] <= 8'hea;
		memory[16'h31cd] <= 8'h1f;
		memory[16'h31ce] <= 8'h2d;
		memory[16'h31cf] <= 8'h95;
		memory[16'h31d0] <= 8'h51;
		memory[16'h31d1] <= 8'h3a;
		memory[16'h31d2] <= 8'hf1;
		memory[16'h31d3] <= 8'h76;
		memory[16'h31d4] <= 8'h65;
		memory[16'h31d5] <= 8'h5;
		memory[16'h31d6] <= 8'h89;
		memory[16'h31d7] <= 8'h2e;
		memory[16'h31d8] <= 8'hdc;
		memory[16'h31d9] <= 8'h23;
		memory[16'h31da] <= 8'hef;
		memory[16'h31db] <= 8'h9;
		memory[16'h31dc] <= 8'h29;
		memory[16'h31dd] <= 8'h2f;
		memory[16'h31de] <= 8'hc6;
		memory[16'h31df] <= 8'h6e;
		memory[16'h31e0] <= 8'hb3;
		memory[16'h31e1] <= 8'ha7;
		memory[16'h31e2] <= 8'hf3;
		memory[16'h31e3] <= 8'h3a;
		memory[16'h31e4] <= 8'h3d;
		memory[16'h31e5] <= 8'he9;
		memory[16'h31e6] <= 8'hd3;
		memory[16'h31e7] <= 8'h33;
		memory[16'h31e8] <= 8'hd5;
		memory[16'h31e9] <= 8'he1;
		memory[16'h31ea] <= 8'h9f;
		memory[16'h31eb] <= 8'hbf;
		memory[16'h31ec] <= 8'h0;
		memory[16'h31ed] <= 8'hcd;
		memory[16'h31ee] <= 8'h55;
		memory[16'h31ef] <= 8'h51;
		memory[16'h31f0] <= 8'h7;
		memory[16'h31f1] <= 8'h46;
		memory[16'h31f2] <= 8'hc8;
		memory[16'h31f3] <= 8'h6d;
		memory[16'h31f4] <= 8'h4b;
		memory[16'h31f5] <= 8'h51;
		memory[16'h31f6] <= 8'h9b;
		memory[16'h31f7] <= 8'h27;
		memory[16'h31f8] <= 8'h74;
		memory[16'h31f9] <= 8'h8a;
		memory[16'h31fa] <= 8'h31;
		memory[16'h31fb] <= 8'h9d;
		memory[16'h31fc] <= 8'hb9;
		memory[16'h31fd] <= 8'hf7;
		memory[16'h31fe] <= 8'hb;
		memory[16'h31ff] <= 8'h6d;
		memory[16'h3200] <= 8'h9f;
		memory[16'h3201] <= 8'hfe;
		memory[16'h3202] <= 8'ha7;
		memory[16'h3203] <= 8'hdc;
		memory[16'h3204] <= 8'he7;
		memory[16'h3205] <= 8'h7b;
		memory[16'h3206] <= 8'hf;
		memory[16'h3207] <= 8'hbd;
		memory[16'h3208] <= 8'h5c;
		memory[16'h3209] <= 8'haf;
		memory[16'h320a] <= 8'h7c;
		memory[16'h320b] <= 8'h5c;
		memory[16'h320c] <= 8'h7c;
		memory[16'h320d] <= 8'hd1;
		memory[16'h320e] <= 8'had;
		memory[16'h320f] <= 8'h83;
		memory[16'h3210] <= 8'h17;
		memory[16'h3211] <= 8'h75;
		memory[16'h3212] <= 8'hf0;
		memory[16'h3213] <= 8'h63;
		memory[16'h3214] <= 8'hc6;
		memory[16'h3215] <= 8'h8b;
		memory[16'h3216] <= 8'h8a;
		memory[16'h3217] <= 8'h3a;
		memory[16'h3218] <= 8'h16;
		memory[16'h3219] <= 8'hbb;
		memory[16'h321a] <= 8'hd7;
		memory[16'h321b] <= 8'hcf;
		memory[16'h321c] <= 8'hb3;
		memory[16'h321d] <= 8'he3;
		memory[16'h321e] <= 8'h3c;
		memory[16'h321f] <= 8'h52;
		memory[16'h3220] <= 8'he1;
		memory[16'h3221] <= 8'he4;
		memory[16'h3222] <= 8'h2e;
		memory[16'h3223] <= 8'hc9;
		memory[16'h3224] <= 8'h5f;
		memory[16'h3225] <= 8'h3e;
		memory[16'h3226] <= 8'h86;
		memory[16'h3227] <= 8'hbb;
		memory[16'h3228] <= 8'hed;
		memory[16'h3229] <= 8'h2;
		memory[16'h322a] <= 8'h17;
		memory[16'h322b] <= 8'h69;
		memory[16'h322c] <= 8'hd4;
		memory[16'h322d] <= 8'hc4;
		memory[16'h322e] <= 8'hec;
		memory[16'h322f] <= 8'heb;
		memory[16'h3230] <= 8'h3a;
		memory[16'h3231] <= 8'hdd;
		memory[16'h3232] <= 8'h4e;
		memory[16'h3233] <= 8'h0;
		memory[16'h3234] <= 8'h68;
		memory[16'h3235] <= 8'hd9;
		memory[16'h3236] <= 8'h3b;
		memory[16'h3237] <= 8'h7e;
		memory[16'h3238] <= 8'h94;
		memory[16'h3239] <= 8'h12;
		memory[16'h323a] <= 8'h4e;
		memory[16'h323b] <= 8'h47;
		memory[16'h323c] <= 8'hf5;
		memory[16'h323d] <= 8'h8a;
		memory[16'h323e] <= 8'h99;
		memory[16'h323f] <= 8'hd7;
		memory[16'h3240] <= 8'h6e;
		memory[16'h3241] <= 8'hc8;
		memory[16'h3242] <= 8'ha0;
		memory[16'h3243] <= 8'hcd;
		memory[16'h3244] <= 8'h6;
		memory[16'h3245] <= 8'h26;
		memory[16'h3246] <= 8'h88;
		memory[16'h3247] <= 8'hf3;
		memory[16'h3248] <= 8'h28;
		memory[16'h3249] <= 8'h9f;
		memory[16'h324a] <= 8'h5c;
		memory[16'h324b] <= 8'hfc;
		memory[16'h324c] <= 8'h64;
		memory[16'h324d] <= 8'h48;
		memory[16'h324e] <= 8'he8;
		memory[16'h324f] <= 8'h9e;
		memory[16'h3250] <= 8'h25;
		memory[16'h3251] <= 8'h36;
		memory[16'h3252] <= 8'h9e;
		memory[16'h3253] <= 8'h8e;
		memory[16'h3254] <= 8'hf;
		memory[16'h3255] <= 8'hd9;
		memory[16'h3256] <= 8'hc;
		memory[16'h3257] <= 8'ha4;
		memory[16'h3258] <= 8'hec;
		memory[16'h3259] <= 8'h5a;
		memory[16'h325a] <= 8'heb;
		memory[16'h325b] <= 8'he1;
		memory[16'h325c] <= 8'he5;
		memory[16'h325d] <= 8'h85;
		memory[16'h325e] <= 8'hb8;
		memory[16'h325f] <= 8'h53;
		memory[16'h3260] <= 8'h4d;
		memory[16'h3261] <= 8'h58;
		memory[16'h3262] <= 8'h21;
		memory[16'h3263] <= 8'h53;
		memory[16'h3264] <= 8'h7e;
		memory[16'h3265] <= 8'ha9;
		memory[16'h3266] <= 8'h46;
		memory[16'h3267] <= 8'ha7;
		memory[16'h3268] <= 8'h49;
		memory[16'h3269] <= 8'ha2;
		memory[16'h326a] <= 8'ha3;
		memory[16'h326b] <= 8'had;
		memory[16'h326c] <= 8'hea;
		memory[16'h326d] <= 8'h8b;
		memory[16'h326e] <= 8'h4b;
		memory[16'h326f] <= 8'h10;
		memory[16'h3270] <= 8'hc2;
		memory[16'h3271] <= 8'he9;
		memory[16'h3272] <= 8'h9e;
		memory[16'h3273] <= 8'hd1;
		memory[16'h3274] <= 8'hc3;
		memory[16'h3275] <= 8'haa;
		memory[16'h3276] <= 8'h75;
		memory[16'h3277] <= 8'haf;
		memory[16'h3278] <= 8'h5;
		memory[16'h3279] <= 8'h61;
		memory[16'h327a] <= 8'h90;
		memory[16'h327b] <= 8'hea;
		memory[16'h327c] <= 8'he6;
		memory[16'h327d] <= 8'h49;
		memory[16'h327e] <= 8'h3d;
		memory[16'h327f] <= 8'h33;
		memory[16'h3280] <= 8'ha1;
		memory[16'h3281] <= 8'h5e;
		memory[16'h3282] <= 8'h86;
		memory[16'h3283] <= 8'h20;
		memory[16'h3284] <= 8'h8;
		memory[16'h3285] <= 8'hcc;
		memory[16'h3286] <= 8'hc7;
		memory[16'h3287] <= 8'h51;
		memory[16'h3288] <= 8'h6e;
		memory[16'h3289] <= 8'h6a;
		memory[16'h328a] <= 8'hfe;
		memory[16'h328b] <= 8'h58;
		memory[16'h328c] <= 8'hf6;
		memory[16'h328d] <= 8'h49;
		memory[16'h328e] <= 8'h68;
		memory[16'h328f] <= 8'hb8;
		memory[16'h3290] <= 8'h32;
		memory[16'h3291] <= 8'h6;
		memory[16'h3292] <= 8'h89;
		memory[16'h3293] <= 8'hf5;
		memory[16'h3294] <= 8'hb1;
		memory[16'h3295] <= 8'hff;
		memory[16'h3296] <= 8'ha4;
		memory[16'h3297] <= 8'hb6;
		memory[16'h3298] <= 8'h60;
		memory[16'h3299] <= 8'h35;
		memory[16'h329a] <= 8'ha0;
		memory[16'h329b] <= 8'h46;
		memory[16'h329c] <= 8'h7e;
		memory[16'h329d] <= 8'hdd;
		memory[16'h329e] <= 8'h79;
		memory[16'h329f] <= 8'h1f;
		memory[16'h32a0] <= 8'h3c;
		memory[16'h32a1] <= 8'hff;
		memory[16'h32a2] <= 8'h3f;
		memory[16'h32a3] <= 8'h44;
		memory[16'h32a4] <= 8'hcb;
		memory[16'h32a5] <= 8'h6;
		memory[16'h32a6] <= 8'h95;
		memory[16'h32a7] <= 8'h39;
		memory[16'h32a8] <= 8'h71;
		memory[16'h32a9] <= 8'h93;
		memory[16'h32aa] <= 8'h91;
		memory[16'h32ab] <= 8'h67;
		memory[16'h32ac] <= 8'hdc;
		memory[16'h32ad] <= 8'hfa;
		memory[16'h32ae] <= 8'h1f;
		memory[16'h32af] <= 8'he;
		memory[16'h32b0] <= 8'h0;
		memory[16'h32b1] <= 8'ha8;
		memory[16'h32b2] <= 8'h4;
		memory[16'h32b3] <= 8'hb1;
		memory[16'h32b4] <= 8'ha7;
		memory[16'h32b5] <= 8'ha8;
		memory[16'h32b6] <= 8'h67;
		memory[16'h32b7] <= 8'h7;
		memory[16'h32b8] <= 8'hdd;
		memory[16'h32b9] <= 8'h7;
		memory[16'h32ba] <= 8'h4d;
		memory[16'h32bb] <= 8'h5b;
		memory[16'h32bc] <= 8'he5;
		memory[16'h32bd] <= 8'hc6;
		memory[16'h32be] <= 8'h7b;
		memory[16'h32bf] <= 8'h21;
		memory[16'h32c0] <= 8'hc5;
		memory[16'h32c1] <= 8'hba;
		memory[16'h32c2] <= 8'h65;
		memory[16'h32c3] <= 8'h90;
		memory[16'h32c4] <= 8'hc1;
		memory[16'h32c5] <= 8'hfa;
		memory[16'h32c6] <= 8'hc9;
		memory[16'h32c7] <= 8'h32;
		memory[16'h32c8] <= 8'h8d;
		memory[16'h32c9] <= 8'h5b;
		memory[16'h32ca] <= 8'h99;
		memory[16'h32cb] <= 8'h69;
		memory[16'h32cc] <= 8'h55;
		memory[16'h32cd] <= 8'hb8;
		memory[16'h32ce] <= 8'h77;
		memory[16'h32cf] <= 8'h55;
		memory[16'h32d0] <= 8'h60;
		memory[16'h32d1] <= 8'h7b;
		memory[16'h32d2] <= 8'h7;
		memory[16'h32d3] <= 8'h8;
		memory[16'h32d4] <= 8'h24;
		memory[16'h32d5] <= 8'h6e;
		memory[16'h32d6] <= 8'hf;
		memory[16'h32d7] <= 8'h1;
		memory[16'h32d8] <= 8'h76;
		memory[16'h32d9] <= 8'h5d;
		memory[16'h32da] <= 8'h5d;
		memory[16'h32db] <= 8'h5b;
		memory[16'h32dc] <= 8'h23;
		memory[16'h32dd] <= 8'hd8;
		memory[16'h32de] <= 8'h7c;
		memory[16'h32df] <= 8'he9;
		memory[16'h32e0] <= 8'h92;
		memory[16'h32e1] <= 8'he1;
		memory[16'h32e2] <= 8'h79;
		memory[16'h32e3] <= 8'h53;
		memory[16'h32e4] <= 8'hdb;
		memory[16'h32e5] <= 8'h43;
		memory[16'h32e6] <= 8'h85;
		memory[16'h32e7] <= 8'h68;
		memory[16'h32e8] <= 8'h9e;
		memory[16'h32e9] <= 8'h1e;
		memory[16'h32ea] <= 8'hd1;
		memory[16'h32eb] <= 8'hf3;
		memory[16'h32ec] <= 8'hd6;
		memory[16'h32ed] <= 8'h48;
		memory[16'h32ee] <= 8'h48;
		memory[16'h32ef] <= 8'h37;
		memory[16'h32f0] <= 8'hc4;
		memory[16'h32f1] <= 8'h4f;
		memory[16'h32f2] <= 8'h3f;
		memory[16'h32f3] <= 8'he8;
		memory[16'h32f4] <= 8'hbe;
		memory[16'h32f5] <= 8'h4e;
		memory[16'h32f6] <= 8'he9;
		memory[16'h32f7] <= 8'h34;
		memory[16'h32f8] <= 8'hab;
		memory[16'h32f9] <= 8'h46;
		memory[16'h32fa] <= 8'h8f;
		memory[16'h32fb] <= 8'hcf;
		memory[16'h32fc] <= 8'h1e;
		memory[16'h32fd] <= 8'hb;
		memory[16'h32fe] <= 8'hb8;
		memory[16'h32ff] <= 8'hb1;
		memory[16'h3300] <= 8'hec;
		memory[16'h3301] <= 8'h31;
		memory[16'h3302] <= 8'h4;
		memory[16'h3303] <= 8'hc7;
		memory[16'h3304] <= 8'h74;
		memory[16'h3305] <= 8'h8a;
		memory[16'h3306] <= 8'h2f;
		memory[16'h3307] <= 8'h12;
		memory[16'h3308] <= 8'ha8;
		memory[16'h3309] <= 8'h0;
		memory[16'h330a] <= 8'h5;
		memory[16'h330b] <= 8'h7f;
		memory[16'h330c] <= 8'h48;
		memory[16'h330d] <= 8'h4e;
		memory[16'h330e] <= 8'hb6;
		memory[16'h330f] <= 8'hc;
		memory[16'h3310] <= 8'h9d;
		memory[16'h3311] <= 8'hf5;
		memory[16'h3312] <= 8'hf4;
		memory[16'h3313] <= 8'h5b;
		memory[16'h3314] <= 8'h43;
		memory[16'h3315] <= 8'hde;
		memory[16'h3316] <= 8'h8f;
		memory[16'h3317] <= 8'hef;
		memory[16'h3318] <= 8'h24;
		memory[16'h3319] <= 8'h1e;
		memory[16'h331a] <= 8'hbe;
		memory[16'h331b] <= 8'h43;
		memory[16'h331c] <= 8'h29;
		memory[16'h331d] <= 8'h76;
		memory[16'h331e] <= 8'hf4;
		memory[16'h331f] <= 8'h15;
		memory[16'h3320] <= 8'ha7;
		memory[16'h3321] <= 8'hf8;
		memory[16'h3322] <= 8'hdc;
		memory[16'h3323] <= 8'h1c;
		memory[16'h3324] <= 8'h82;
		memory[16'h3325] <= 8'hb;
		memory[16'h3326] <= 8'h2e;
		memory[16'h3327] <= 8'h2b;
		memory[16'h3328] <= 8'hb;
		memory[16'h3329] <= 8'h34;
		memory[16'h332a] <= 8'haa;
		memory[16'h332b] <= 8'h54;
		memory[16'h332c] <= 8'h82;
		memory[16'h332d] <= 8'h60;
		memory[16'h332e] <= 8'h60;
		memory[16'h332f] <= 8'h1f;
		memory[16'h3330] <= 8'h55;
		memory[16'h3331] <= 8'h55;
		memory[16'h3332] <= 8'h7b;
		memory[16'h3333] <= 8'h98;
		memory[16'h3334] <= 8'h33;
		memory[16'h3335] <= 8'ha;
		memory[16'h3336] <= 8'h87;
		memory[16'h3337] <= 8'h57;
		memory[16'h3338] <= 8'h29;
		memory[16'h3339] <= 8'h45;
		memory[16'h333a] <= 8'h9a;
		memory[16'h333b] <= 8'h52;
		memory[16'h333c] <= 8'hbb;
		memory[16'h333d] <= 8'h8e;
		memory[16'h333e] <= 8'h68;
		memory[16'h333f] <= 8'h63;
		memory[16'h3340] <= 8'h87;
		memory[16'h3341] <= 8'h44;
		memory[16'h3342] <= 8'h7f;
		memory[16'h3343] <= 8'h9;
		memory[16'h3344] <= 8'h50;
		memory[16'h3345] <= 8'had;
		memory[16'h3346] <= 8'h34;
		memory[16'h3347] <= 8'h5b;
		memory[16'h3348] <= 8'he1;
		memory[16'h3349] <= 8'hde;
		memory[16'h334a] <= 8'haf;
		memory[16'h334b] <= 8'h63;
		memory[16'h334c] <= 8'h3e;
		memory[16'h334d] <= 8'h10;
		memory[16'h334e] <= 8'h83;
		memory[16'h334f] <= 8'h93;
		memory[16'h3350] <= 8'h65;
		memory[16'h3351] <= 8'hfe;
		memory[16'h3352] <= 8'h2c;
		memory[16'h3353] <= 8'h98;
		memory[16'h3354] <= 8'h8;
		memory[16'h3355] <= 8'hb3;
		memory[16'h3356] <= 8'hef;
		memory[16'h3357] <= 8'h31;
		memory[16'h3358] <= 8'hf9;
		memory[16'h3359] <= 8'h8a;
		memory[16'h335a] <= 8'h84;
		memory[16'h335b] <= 8'hb4;
		memory[16'h335c] <= 8'h18;
		memory[16'h335d] <= 8'hec;
		memory[16'h335e] <= 8'h17;
		memory[16'h335f] <= 8'h9f;
		memory[16'h3360] <= 8'h30;
		memory[16'h3361] <= 8'h96;
		memory[16'h3362] <= 8'ha9;
		memory[16'h3363] <= 8'h80;
		memory[16'h3364] <= 8'h44;
		memory[16'h3365] <= 8'hdd;
		memory[16'h3366] <= 8'hdc;
		memory[16'h3367] <= 8'h25;
		memory[16'h3368] <= 8'hbc;
		memory[16'h3369] <= 8'h8b;
		memory[16'h336a] <= 8'h89;
		memory[16'h336b] <= 8'hfa;
		memory[16'h336c] <= 8'h9b;
		memory[16'h336d] <= 8'hc;
		memory[16'h336e] <= 8'h8e;
		memory[16'h336f] <= 8'h0;
		memory[16'h3370] <= 8'ha;
		memory[16'h3371] <= 8'hba;
		memory[16'h3372] <= 8'h98;
		memory[16'h3373] <= 8'h12;
		memory[16'h3374] <= 8'h6d;
		memory[16'h3375] <= 8'h88;
		memory[16'h3376] <= 8'h44;
		memory[16'h3377] <= 8'h66;
		memory[16'h3378] <= 8'h12;
		memory[16'h3379] <= 8'hc8;
		memory[16'h337a] <= 8'h1b;
		memory[16'h337b] <= 8'h2a;
		memory[16'h337c] <= 8'hb4;
		memory[16'h337d] <= 8'h32;
		memory[16'h337e] <= 8'hca;
		memory[16'h337f] <= 8'he4;
		memory[16'h3380] <= 8'hc9;
		memory[16'h3381] <= 8'h73;
		memory[16'h3382] <= 8'h65;
		memory[16'h3383] <= 8'hd;
		memory[16'h3384] <= 8'h50;
		memory[16'h3385] <= 8'h41;
		memory[16'h3386] <= 8'h32;
		memory[16'h3387] <= 8'hc;
		memory[16'h3388] <= 8'hcc;
		memory[16'h3389] <= 8'hbb;
		memory[16'h338a] <= 8'h7;
		memory[16'h338b] <= 8'h68;
		memory[16'h338c] <= 8'hc7;
		memory[16'h338d] <= 8'h95;
		memory[16'h338e] <= 8'h68;
		memory[16'h338f] <= 8'hd1;
		memory[16'h3390] <= 8'h4f;
		memory[16'h3391] <= 8'h1;
		memory[16'h3392] <= 8'he4;
		memory[16'h3393] <= 8'hbc;
		memory[16'h3394] <= 8'h89;
		memory[16'h3395] <= 8'h28;
		memory[16'h3396] <= 8'h23;
		memory[16'h3397] <= 8'h9b;
		memory[16'h3398] <= 8'hf0;
		memory[16'h3399] <= 8'h3e;
		memory[16'h339a] <= 8'hc5;
		memory[16'h339b] <= 8'ha4;
		memory[16'h339c] <= 8'h70;
		memory[16'h339d] <= 8'h8f;
		memory[16'h339e] <= 8'h88;
		memory[16'h339f] <= 8'h39;
		memory[16'h33a0] <= 8'h2;
		memory[16'h33a1] <= 8'hed;
		memory[16'h33a2] <= 8'h46;
		memory[16'h33a3] <= 8'h53;
		memory[16'h33a4] <= 8'h2e;
		memory[16'h33a5] <= 8'h79;
		memory[16'h33a6] <= 8'h5f;
		memory[16'h33a7] <= 8'hfb;
		memory[16'h33a8] <= 8'h34;
		memory[16'h33a9] <= 8'h66;
		memory[16'h33aa] <= 8'h63;
		memory[16'h33ab] <= 8'hfc;
		memory[16'h33ac] <= 8'hfb;
		memory[16'h33ad] <= 8'hcb;
		memory[16'h33ae] <= 8'hcd;
		memory[16'h33af] <= 8'h4a;
		memory[16'h33b0] <= 8'hcc;
		memory[16'h33b1] <= 8'hb1;
		memory[16'h33b2] <= 8'h7;
		memory[16'h33b3] <= 8'h55;
		memory[16'h33b4] <= 8'hd9;
		memory[16'h33b5] <= 8'h2a;
		memory[16'h33b6] <= 8'hf0;
		memory[16'h33b7] <= 8'hc9;
		memory[16'h33b8] <= 8'h68;
		memory[16'h33b9] <= 8'hb6;
		memory[16'h33ba] <= 8'h6d;
		memory[16'h33bb] <= 8'hd8;
		memory[16'h33bc] <= 8'h45;
		memory[16'h33bd] <= 8'hf6;
		memory[16'h33be] <= 8'h12;
		memory[16'h33bf] <= 8'h48;
		memory[16'h33c0] <= 8'he3;
		memory[16'h33c1] <= 8'h58;
		memory[16'h33c2] <= 8'h9b;
		memory[16'h33c3] <= 8'h12;
		memory[16'h33c4] <= 8'hd1;
		memory[16'h33c5] <= 8'hfa;
		memory[16'h33c6] <= 8'hd;
		memory[16'h33c7] <= 8'h6;
		memory[16'h33c8] <= 8'h61;
		memory[16'h33c9] <= 8'h70;
		memory[16'h33ca] <= 8'h2;
		memory[16'h33cb] <= 8'h5c;
		memory[16'h33cc] <= 8'h3b;
		memory[16'h33cd] <= 8'hcf;
		memory[16'h33ce] <= 8'ha7;
		memory[16'h33cf] <= 8'h8;
		memory[16'h33d0] <= 8'h81;
		memory[16'h33d1] <= 8'hae;
		memory[16'h33d2] <= 8'h5d;
		memory[16'h33d3] <= 8'h5a;
		memory[16'h33d4] <= 8'hd8;
		memory[16'h33d5] <= 8'h4e;
		memory[16'h33d6] <= 8'h24;
		memory[16'h33d7] <= 8'h40;
		memory[16'h33d8] <= 8'h4;
		memory[16'h33d9] <= 8'h91;
		memory[16'h33da] <= 8'h18;
		memory[16'h33db] <= 8'h49;
		memory[16'h33dc] <= 8'h87;
		memory[16'h33dd] <= 8'h2a;
		memory[16'h33de] <= 8'h91;
		memory[16'h33df] <= 8'h6b;
		memory[16'h33e0] <= 8'h83;
		memory[16'h33e1] <= 8'h2c;
		memory[16'h33e2] <= 8'h7d;
		memory[16'h33e3] <= 8'h54;
		memory[16'h33e4] <= 8'h27;
		memory[16'h33e5] <= 8'h8a;
		memory[16'h33e6] <= 8'h5a;
		memory[16'h33e7] <= 8'h88;
		memory[16'h33e8] <= 8'hfa;
		memory[16'h33e9] <= 8'h5c;
		memory[16'h33ea] <= 8'he4;
		memory[16'h33eb] <= 8'h35;
		memory[16'h33ec] <= 8'h2c;
		memory[16'h33ed] <= 8'h8b;
		memory[16'h33ee] <= 8'h3d;
		memory[16'h33ef] <= 8'had;
		memory[16'h33f0] <= 8'h39;
		memory[16'h33f1] <= 8'h9b;
		memory[16'h33f2] <= 8'h7;
		memory[16'h33f3] <= 8'h11;
		memory[16'h33f4] <= 8'he9;
		memory[16'h33f5] <= 8'h2b;
		memory[16'h33f6] <= 8'h51;
		memory[16'h33f7] <= 8'hed;
		memory[16'h33f8] <= 8'hbd;
		memory[16'h33f9] <= 8'h6a;
		memory[16'h33fa] <= 8'h36;
		memory[16'h33fb] <= 8'h44;
		memory[16'h33fc] <= 8'h94;
		memory[16'h33fd] <= 8'hc8;
		memory[16'h33fe] <= 8'haf;
		memory[16'h33ff] <= 8'h17;
		memory[16'h3400] <= 8'hf4;
		memory[16'h3401] <= 8'h2c;
		memory[16'h3402] <= 8'h6c;
		memory[16'h3403] <= 8'h1b;
		memory[16'h3404] <= 8'hb6;
		memory[16'h3405] <= 8'hc6;
		memory[16'h3406] <= 8'ha3;
		memory[16'h3407] <= 8'hb0;
		memory[16'h3408] <= 8'h23;
		memory[16'h3409] <= 8'h88;
		memory[16'h340a] <= 8'he6;
		memory[16'h340b] <= 8'h4f;
		memory[16'h340c] <= 8'h13;
		memory[16'h340d] <= 8'h23;
		memory[16'h340e] <= 8'hfc;
		memory[16'h340f] <= 8'h4d;
		memory[16'h3410] <= 8'hbe;
		memory[16'h3411] <= 8'h3;
		memory[16'h3412] <= 8'h5e;
		memory[16'h3413] <= 8'ha7;
		memory[16'h3414] <= 8'h2f;
		memory[16'h3415] <= 8'hb0;
		memory[16'h3416] <= 8'h94;
		memory[16'h3417] <= 8'hec;
		memory[16'h3418] <= 8'h1a;
		memory[16'h3419] <= 8'hcb;
		memory[16'h341a] <= 8'h30;
		memory[16'h341b] <= 8'hae;
		memory[16'h341c] <= 8'h93;
		memory[16'h341d] <= 8'he0;
		memory[16'h341e] <= 8'hc6;
		memory[16'h341f] <= 8'h87;
		memory[16'h3420] <= 8'hc;
		memory[16'h3421] <= 8'h32;
		memory[16'h3422] <= 8'ha3;
		memory[16'h3423] <= 8'hc3;
		memory[16'h3424] <= 8'hf8;
		memory[16'h3425] <= 8'h46;
		memory[16'h3426] <= 8'h73;
		memory[16'h3427] <= 8'h1b;
		memory[16'h3428] <= 8'hce;
		memory[16'h3429] <= 8'h59;
		memory[16'h342a] <= 8'h6a;
		memory[16'h342b] <= 8'he2;
		memory[16'h342c] <= 8'h7d;
		memory[16'h342d] <= 8'h66;
		memory[16'h342e] <= 8'h2f;
		memory[16'h342f] <= 8'h3b;
		memory[16'h3430] <= 8'h6a;
		memory[16'h3431] <= 8'h8d;
		memory[16'h3432] <= 8'he3;
		memory[16'h3433] <= 8'h99;
		memory[16'h3434] <= 8'h3d;
		memory[16'h3435] <= 8'h77;
		memory[16'h3436] <= 8'h85;
		memory[16'h3437] <= 8'h57;
		memory[16'h3438] <= 8'h42;
		memory[16'h3439] <= 8'hb5;
		memory[16'h343a] <= 8'h6;
		memory[16'h343b] <= 8'hd5;
		memory[16'h343c] <= 8'h95;
		memory[16'h343d] <= 8'hcc;
		memory[16'h343e] <= 8'h5d;
		memory[16'h343f] <= 8'ha2;
		memory[16'h3440] <= 8'hfe;
		memory[16'h3441] <= 8'h0;
		memory[16'h3442] <= 8'h65;
		memory[16'h3443] <= 8'hf6;
		memory[16'h3444] <= 8'h46;
		memory[16'h3445] <= 8'hd8;
		memory[16'h3446] <= 8'h12;
		memory[16'h3447] <= 8'h15;
		memory[16'h3448] <= 8'h32;
		memory[16'h3449] <= 8'h7c;
		memory[16'h344a] <= 8'hf7;
		memory[16'h344b] <= 8'haf;
		memory[16'h344c] <= 8'he3;
		memory[16'h344d] <= 8'h26;
		memory[16'h344e] <= 8'hea;
		memory[16'h344f] <= 8'h4d;
		memory[16'h3450] <= 8'hb3;
		memory[16'h3451] <= 8'hcd;
		memory[16'h3452] <= 8'he6;
		memory[16'h3453] <= 8'hf1;
		memory[16'h3454] <= 8'h45;
		memory[16'h3455] <= 8'h6b;
		memory[16'h3456] <= 8'h48;
		memory[16'h3457] <= 8'h87;
		memory[16'h3458] <= 8'h20;
		memory[16'h3459] <= 8'h4e;
		memory[16'h345a] <= 8'h5d;
		memory[16'h345b] <= 8'hb6;
		memory[16'h345c] <= 8'h1a;
		memory[16'h345d] <= 8'hba;
		memory[16'h345e] <= 8'h58;
		memory[16'h345f] <= 8'h18;
		memory[16'h3460] <= 8'hba;
		memory[16'h3461] <= 8'hbd;
		memory[16'h3462] <= 8'hf;
		memory[16'h3463] <= 8'h0;
		memory[16'h3464] <= 8'h95;
		memory[16'h3465] <= 8'h21;
		memory[16'h3466] <= 8'h15;
		memory[16'h3467] <= 8'hc7;
		memory[16'h3468] <= 8'h9d;
		memory[16'h3469] <= 8'hc;
		memory[16'h346a] <= 8'h76;
		memory[16'h346b] <= 8'h80;
		memory[16'h346c] <= 8'h32;
		memory[16'h346d] <= 8'h61;
		memory[16'h346e] <= 8'hcd;
		memory[16'h346f] <= 8'he6;
		memory[16'h3470] <= 8'h2e;
		memory[16'h3471] <= 8'hb3;
		memory[16'h3472] <= 8'hd7;
		memory[16'h3473] <= 8'h73;
		memory[16'h3474] <= 8'h1e;
		memory[16'h3475] <= 8'h1f;
		memory[16'h3476] <= 8'hfb;
		memory[16'h3477] <= 8'h3f;
		memory[16'h3478] <= 8'h6e;
		memory[16'h3479] <= 8'h58;
		memory[16'h347a] <= 8'hf5;
		memory[16'h347b] <= 8'h88;
		memory[16'h347c] <= 8'h12;
		memory[16'h347d] <= 8'h4d;
		memory[16'h347e] <= 8'ha1;
		memory[16'h347f] <= 8'hcc;
		memory[16'h3480] <= 8'ha;
		memory[16'h3481] <= 8'hb0;
		memory[16'h3482] <= 8'hcc;
		memory[16'h3483] <= 8'h9f;
		memory[16'h3484] <= 8'hd1;
		memory[16'h3485] <= 8'he2;
		memory[16'h3486] <= 8'h67;
		memory[16'h3487] <= 8'h6e;
		memory[16'h3488] <= 8'hee;
		memory[16'h3489] <= 8'hdd;
		memory[16'h348a] <= 8'hef;
		memory[16'h348b] <= 8'h21;
		memory[16'h348c] <= 8'h3e;
		memory[16'h348d] <= 8'hbc;
		memory[16'h348e] <= 8'h7;
		memory[16'h348f] <= 8'h6d;
		memory[16'h3490] <= 8'h70;
		memory[16'h3491] <= 8'hde;
		memory[16'h3492] <= 8'he0;
		memory[16'h3493] <= 8'h8e;
		memory[16'h3494] <= 8'hfd;
		memory[16'h3495] <= 8'hdb;
		memory[16'h3496] <= 8'hcd;
		memory[16'h3497] <= 8'h6b;
		memory[16'h3498] <= 8'h33;
		memory[16'h3499] <= 8'hc2;
		memory[16'h349a] <= 8'hf4;
		memory[16'h349b] <= 8'h45;
		memory[16'h349c] <= 8'hf;
		memory[16'h349d] <= 8'h95;
		memory[16'h349e] <= 8'h11;
		memory[16'h349f] <= 8'h19;
		memory[16'h34a0] <= 8'h45;
		memory[16'h34a1] <= 8'hde;
		memory[16'h34a2] <= 8'hb9;
		memory[16'h34a3] <= 8'h16;
		memory[16'h34a4] <= 8'hc0;
		memory[16'h34a5] <= 8'h20;
		memory[16'h34a6] <= 8'h84;
		memory[16'h34a7] <= 8'hae;
		memory[16'h34a8] <= 8'hfd;
		memory[16'h34a9] <= 8'h73;
		memory[16'h34aa] <= 8'hcf;
		memory[16'h34ab] <= 8'h3c;
		memory[16'h34ac] <= 8'h30;
		memory[16'h34ad] <= 8'hd6;
		memory[16'h34ae] <= 8'ha9;
		memory[16'h34af] <= 8'ha0;
		memory[16'h34b0] <= 8'hb4;
		memory[16'h34b1] <= 8'h89;
		memory[16'h34b2] <= 8'h2e;
		memory[16'h34b3] <= 8'hb2;
		memory[16'h34b4] <= 8'h65;
		memory[16'h34b5] <= 8'hfc;
		memory[16'h34b6] <= 8'h1d;
		memory[16'h34b7] <= 8'h98;
		memory[16'h34b8] <= 8'hbe;
		memory[16'h34b9] <= 8'h11;
		memory[16'h34ba] <= 8'hde;
		memory[16'h34bb] <= 8'hce;
		memory[16'h34bc] <= 8'ha6;
		memory[16'h34bd] <= 8'hef;
		memory[16'h34be] <= 8'he7;
		memory[16'h34bf] <= 8'heb;
		memory[16'h34c0] <= 8'hcd;
		memory[16'h34c1] <= 8'ha0;
		memory[16'h34c2] <= 8'h1;
		memory[16'h34c3] <= 8'h8d;
		memory[16'h34c4] <= 8'hc0;
		memory[16'h34c5] <= 8'h86;
		memory[16'h34c6] <= 8'h3c;
		memory[16'h34c7] <= 8'hbe;
		memory[16'h34c8] <= 8'hf9;
		memory[16'h34c9] <= 8'hb;
		memory[16'h34ca] <= 8'hfa;
		memory[16'h34cb] <= 8'h29;
		memory[16'h34cc] <= 8'he2;
		memory[16'h34cd] <= 8'ha3;
		memory[16'h34ce] <= 8'hc9;
		memory[16'h34cf] <= 8'h96;
		memory[16'h34d0] <= 8'h2c;
		memory[16'h34d1] <= 8'hf8;
		memory[16'h34d2] <= 8'h48;
		memory[16'h34d3] <= 8'h91;
		memory[16'h34d4] <= 8'hf4;
		memory[16'h34d5] <= 8'h66;
		memory[16'h34d6] <= 8'h2a;
		memory[16'h34d7] <= 8'hb2;
		memory[16'h34d8] <= 8'h77;
		memory[16'h34d9] <= 8'h8;
		memory[16'h34da] <= 8'h80;
		memory[16'h34db] <= 8'h1e;
		memory[16'h34dc] <= 8'hf7;
		memory[16'h34dd] <= 8'h68;
		memory[16'h34de] <= 8'h9;
		memory[16'h34df] <= 8'hc5;
		memory[16'h34e0] <= 8'h8;
		memory[16'h34e1] <= 8'hb;
		memory[16'h34e2] <= 8'h52;
		memory[16'h34e3] <= 8'hc9;
		memory[16'h34e4] <= 8'h91;
		memory[16'h34e5] <= 8'h8e;
		memory[16'h34e6] <= 8'h87;
		memory[16'h34e7] <= 8'h8a;
		memory[16'h34e8] <= 8'h9a;
		memory[16'h34e9] <= 8'h81;
		memory[16'h34ea] <= 8'hb4;
		memory[16'h34eb] <= 8'h7c;
		memory[16'h34ec] <= 8'h24;
		memory[16'h34ed] <= 8'h7d;
		memory[16'h34ee] <= 8'h12;
		memory[16'h34ef] <= 8'h50;
		memory[16'h34f0] <= 8'h75;
		memory[16'h34f1] <= 8'h5b;
		memory[16'h34f2] <= 8'he2;
		memory[16'h34f3] <= 8'h69;
		memory[16'h34f4] <= 8'hc1;
		memory[16'h34f5] <= 8'hc;
		memory[16'h34f6] <= 8'h1c;
		memory[16'h34f7] <= 8'h38;
		memory[16'h34f8] <= 8'h14;
		memory[16'h34f9] <= 8'h9c;
		memory[16'h34fa] <= 8'h56;
		memory[16'h34fb] <= 8'hb;
		memory[16'h34fc] <= 8'h4;
		memory[16'h34fd] <= 8'h60;
		memory[16'h34fe] <= 8'hd0;
		memory[16'h34ff] <= 8'hd;
		memory[16'h3500] <= 8'h6b;
		memory[16'h3501] <= 8'h23;
		memory[16'h3502] <= 8'hd6;
		memory[16'h3503] <= 8'hfc;
		memory[16'h3504] <= 8'hb1;
		memory[16'h3505] <= 8'h5d;
		memory[16'h3506] <= 8'h86;
		memory[16'h3507] <= 8'h4b;
		memory[16'h3508] <= 8'hde;
		memory[16'h3509] <= 8'h3a;
		memory[16'h350a] <= 8'hc7;
		memory[16'h350b] <= 8'h2;
		memory[16'h350c] <= 8'hb8;
		memory[16'h350d] <= 8'hda;
		memory[16'h350e] <= 8'h52;
		memory[16'h350f] <= 8'h2d;
		memory[16'h3510] <= 8'h35;
		memory[16'h3511] <= 8'h34;
		memory[16'h3512] <= 8'h97;
		memory[16'h3513] <= 8'hf6;
		memory[16'h3514] <= 8'h40;
		memory[16'h3515] <= 8'hb3;
		memory[16'h3516] <= 8'h2e;
		memory[16'h3517] <= 8'h54;
		memory[16'h3518] <= 8'h4f;
		memory[16'h3519] <= 8'h85;
		memory[16'h351a] <= 8'h60;
		memory[16'h351b] <= 8'h54;
		memory[16'h351c] <= 8'he5;
		memory[16'h351d] <= 8'h30;
		memory[16'h351e] <= 8'h61;
		memory[16'h351f] <= 8'h50;
		memory[16'h3520] <= 8'h53;
		memory[16'h3521] <= 8'h37;
		memory[16'h3522] <= 8'h4c;
		memory[16'h3523] <= 8'h5;
		memory[16'h3524] <= 8'h94;
		memory[16'h3525] <= 8'hd2;
		memory[16'h3526] <= 8'h50;
		memory[16'h3527] <= 8'h72;
		memory[16'h3528] <= 8'hd;
		memory[16'h3529] <= 8'h18;
		memory[16'h352a] <= 8'h74;
		memory[16'h352b] <= 8'hc5;
		memory[16'h352c] <= 8'hf2;
		memory[16'h352d] <= 8'hc6;
		memory[16'h352e] <= 8'hf2;
		memory[16'h352f] <= 8'h27;
		memory[16'h3530] <= 8'hfb;
		memory[16'h3531] <= 8'h89;
		memory[16'h3532] <= 8'h1d;
		memory[16'h3533] <= 8'h3b;
		memory[16'h3534] <= 8'h3c;
		memory[16'h3535] <= 8'h4b;
		memory[16'h3536] <= 8'h90;
		memory[16'h3537] <= 8'h8c;
		memory[16'h3538] <= 8'hd0;
		memory[16'h3539] <= 8'hf0;
		memory[16'h353a] <= 8'he0;
		memory[16'h353b] <= 8'hb5;
		memory[16'h353c] <= 8'h20;
		memory[16'h353d] <= 8'h41;
		memory[16'h353e] <= 8'h5;
		memory[16'h353f] <= 8'h74;
		memory[16'h3540] <= 8'h78;
		memory[16'h3541] <= 8'h51;
		memory[16'h3542] <= 8'h79;
		memory[16'h3543] <= 8'hc;
		memory[16'h3544] <= 8'h24;
		memory[16'h3545] <= 8'hc9;
		memory[16'h3546] <= 8'h7e;
		memory[16'h3547] <= 8'h31;
		memory[16'h3548] <= 8'he1;
		memory[16'h3549] <= 8'hf2;
		memory[16'h354a] <= 8'hf6;
		memory[16'h354b] <= 8'hd3;
		memory[16'h354c] <= 8'hb8;
		memory[16'h354d] <= 8'he8;
		memory[16'h354e] <= 8'hfa;
		memory[16'h354f] <= 8'hb3;
		memory[16'h3550] <= 8'h72;
		memory[16'h3551] <= 8'h17;
		memory[16'h3552] <= 8'hef;
		memory[16'h3553] <= 8'hae;
		memory[16'h3554] <= 8'h63;
		memory[16'h3555] <= 8'h7f;
		memory[16'h3556] <= 8'h3a;
		memory[16'h3557] <= 8'h33;
		memory[16'h3558] <= 8'h6f;
		memory[16'h3559] <= 8'h1a;
		memory[16'h355a] <= 8'he9;
		memory[16'h355b] <= 8'h8f;
		memory[16'h355c] <= 8'h5b;
		memory[16'h355d] <= 8'hee;
		memory[16'h355e] <= 8'h3;
		memory[16'h355f] <= 8'hd3;
		memory[16'h3560] <= 8'h40;
		memory[16'h3561] <= 8'h7c;
		memory[16'h3562] <= 8'hdf;
		memory[16'h3563] <= 8'h64;
		memory[16'h3564] <= 8'h46;
		memory[16'h3565] <= 8'h5d;
		memory[16'h3566] <= 8'h95;
		memory[16'h3567] <= 8'h27;
		memory[16'h3568] <= 8'h4f;
		memory[16'h3569] <= 8'h8b;
		memory[16'h356a] <= 8'hfb;
		memory[16'h356b] <= 8'h8;
		memory[16'h356c] <= 8'h73;
		memory[16'h356d] <= 8'hf5;
		memory[16'h356e] <= 8'hbb;
		memory[16'h356f] <= 8'he5;
		memory[16'h3570] <= 8'hd;
		memory[16'h3571] <= 8'haa;
		memory[16'h3572] <= 8'h94;
		memory[16'h3573] <= 8'h70;
		memory[16'h3574] <= 8'h29;
		memory[16'h3575] <= 8'hce;
		memory[16'h3576] <= 8'ha3;
		memory[16'h3577] <= 8'h98;
		memory[16'h3578] <= 8'he9;
		memory[16'h3579] <= 8'h8c;
		memory[16'h357a] <= 8'h28;
		memory[16'h357b] <= 8'h44;
		memory[16'h357c] <= 8'h7b;
		memory[16'h357d] <= 8'h2b;
		memory[16'h357e] <= 8'h18;
		memory[16'h357f] <= 8'hbb;
		memory[16'h3580] <= 8'ha8;
		memory[16'h3581] <= 8'hf7;
		memory[16'h3582] <= 8'h1f;
		memory[16'h3583] <= 8'hee;
		memory[16'h3584] <= 8'h55;
		memory[16'h3585] <= 8'hb4;
		memory[16'h3586] <= 8'h15;
		memory[16'h3587] <= 8'ha4;
		memory[16'h3588] <= 8'h3f;
		memory[16'h3589] <= 8'h10;
		memory[16'h358a] <= 8'hac;
		memory[16'h358b] <= 8'hb2;
		memory[16'h358c] <= 8'h6;
		memory[16'h358d] <= 8'h68;
		memory[16'h358e] <= 8'h98;
		memory[16'h358f] <= 8'h13;
		memory[16'h3590] <= 8'h12;
		memory[16'h3591] <= 8'h2c;
		memory[16'h3592] <= 8'h83;
		memory[16'h3593] <= 8'h3c;
		memory[16'h3594] <= 8'hfa;
		memory[16'h3595] <= 8'h26;
		memory[16'h3596] <= 8'hd4;
		memory[16'h3597] <= 8'he3;
		memory[16'h3598] <= 8'hb3;
		memory[16'h3599] <= 8'hfc;
		memory[16'h359a] <= 8'h28;
		memory[16'h359b] <= 8'h2e;
		memory[16'h359c] <= 8'h28;
		memory[16'h359d] <= 8'h40;
		memory[16'h359e] <= 8'he9;
		memory[16'h359f] <= 8'hd0;
		memory[16'h35a0] <= 8'h37;
		memory[16'h35a1] <= 8'h8;
		memory[16'h35a2] <= 8'hbe;
		memory[16'h35a3] <= 8'h8c;
		memory[16'h35a4] <= 8'hbc;
		memory[16'h35a5] <= 8'hd3;
		memory[16'h35a6] <= 8'h31;
		memory[16'h35a7] <= 8'hfb;
		memory[16'h35a8] <= 8'he4;
		memory[16'h35a9] <= 8'hdd;
		memory[16'h35aa] <= 8'had;
		memory[16'h35ab] <= 8'hea;
		memory[16'h35ac] <= 8'h45;
		memory[16'h35ad] <= 8'h45;
		memory[16'h35ae] <= 8'hfd;
		memory[16'h35af] <= 8'h58;
		memory[16'h35b0] <= 8'h71;
		memory[16'h35b1] <= 8'h80;
		memory[16'h35b2] <= 8'h94;
		memory[16'h35b3] <= 8'h6c;
		memory[16'h35b4] <= 8'ha6;
		memory[16'h35b5] <= 8'h68;
		memory[16'h35b6] <= 8'h4f;
		memory[16'h35b7] <= 8'h59;
		memory[16'h35b8] <= 8'h65;
		memory[16'h35b9] <= 8'h77;
		memory[16'h35ba] <= 8'h87;
		memory[16'h35bb] <= 8'h8d;
		memory[16'h35bc] <= 8'hb7;
		memory[16'h35bd] <= 8'h70;
		memory[16'h35be] <= 8'h5d;
		memory[16'h35bf] <= 8'hef;
		memory[16'h35c0] <= 8'h78;
		memory[16'h35c1] <= 8'h1b;
		memory[16'h35c2] <= 8'h7b;
		memory[16'h35c3] <= 8'h34;
		memory[16'h35c4] <= 8'hee;
		memory[16'h35c5] <= 8'hac;
		memory[16'h35c6] <= 8'h2f;
		memory[16'h35c7] <= 8'hd2;
		memory[16'h35c8] <= 8'h8a;
		memory[16'h35c9] <= 8'hdd;
		memory[16'h35ca] <= 8'hbc;
		memory[16'h35cb] <= 8'hcf;
		memory[16'h35cc] <= 8'h22;
		memory[16'h35cd] <= 8'hb9;
		memory[16'h35ce] <= 8'h27;
		memory[16'h35cf] <= 8'h94;
		memory[16'h35d0] <= 8'h39;
		memory[16'h35d1] <= 8'hbb;
		memory[16'h35d2] <= 8'h0;
		memory[16'h35d3] <= 8'he0;
		memory[16'h35d4] <= 8'h24;
		memory[16'h35d5] <= 8'h4f;
		memory[16'h35d6] <= 8'h39;
		memory[16'h35d7] <= 8'h89;
		memory[16'h35d8] <= 8'hc7;
		memory[16'h35d9] <= 8'hc1;
		memory[16'h35da] <= 8'h16;
		memory[16'h35db] <= 8'h7e;
		memory[16'h35dc] <= 8'h31;
		memory[16'h35dd] <= 8'h73;
		memory[16'h35de] <= 8'h6d;
		memory[16'h35df] <= 8'haa;
		memory[16'h35e0] <= 8'h8e;
		memory[16'h35e1] <= 8'he9;
		memory[16'h35e2] <= 8'hde;
		memory[16'h35e3] <= 8'h7c;
		memory[16'h35e4] <= 8'h95;
		memory[16'h35e5] <= 8'he;
		memory[16'h35e6] <= 8'h4f;
		memory[16'h35e7] <= 8'h1f;
		memory[16'h35e8] <= 8'heb;
		memory[16'h35e9] <= 8'hb;
		memory[16'h35ea] <= 8'hef;
		memory[16'h35eb] <= 8'hd;
		memory[16'h35ec] <= 8'hc5;
		memory[16'h35ed] <= 8'h16;
		memory[16'h35ee] <= 8'ha1;
		memory[16'h35ef] <= 8'hfe;
		memory[16'h35f0] <= 8'hd2;
		memory[16'h35f1] <= 8'ha1;
		memory[16'h35f2] <= 8'hde;
		memory[16'h35f3] <= 8'hf6;
		memory[16'h35f4] <= 8'hf1;
		memory[16'h35f5] <= 8'h18;
		memory[16'h35f6] <= 8'h7f;
		memory[16'h35f7] <= 8'hb8;
		memory[16'h35f8] <= 8'hd9;
		memory[16'h35f9] <= 8'h95;
		memory[16'h35fa] <= 8'h36;
		memory[16'h35fb] <= 8'ha;
		memory[16'h35fc] <= 8'h8;
		memory[16'h35fd] <= 8'ha4;
		memory[16'h35fe] <= 8'hb4;
		memory[16'h35ff] <= 8'h96;
		memory[16'h3600] <= 8'h8d;
		memory[16'h3601] <= 8'h93;
		memory[16'h3602] <= 8'h12;
		memory[16'h3603] <= 8'h22;
		memory[16'h3604] <= 8'ha1;
		memory[16'h3605] <= 8'h61;
		memory[16'h3606] <= 8'h42;
		memory[16'h3607] <= 8'h8c;
		memory[16'h3608] <= 8'h6d;
		memory[16'h3609] <= 8'h31;
		memory[16'h360a] <= 8'h99;
		memory[16'h360b] <= 8'h32;
		memory[16'h360c] <= 8'h47;
		memory[16'h360d] <= 8'h3b;
		memory[16'h360e] <= 8'h30;
		memory[16'h360f] <= 8'h19;
		memory[16'h3610] <= 8'hdc;
		memory[16'h3611] <= 8'hf;
		memory[16'h3612] <= 8'hf;
		memory[16'h3613] <= 8'hcd;
		memory[16'h3614] <= 8'h27;
		memory[16'h3615] <= 8'h8e;
		memory[16'h3616] <= 8'h85;
		memory[16'h3617] <= 8'h0;
		memory[16'h3618] <= 8'h23;
		memory[16'h3619] <= 8'hbc;
		memory[16'h361a] <= 8'ha;
		memory[16'h361b] <= 8'h2b;
		memory[16'h361c] <= 8'h60;
		memory[16'h361d] <= 8'hbf;
		memory[16'h361e] <= 8'hc1;
		memory[16'h361f] <= 8'hed;
		memory[16'h3620] <= 8'h52;
		memory[16'h3621] <= 8'hd4;
		memory[16'h3622] <= 8'hf;
		memory[16'h3623] <= 8'hf3;
		memory[16'h3624] <= 8'h35;
		memory[16'h3625] <= 8'h51;
		memory[16'h3626] <= 8'h7f;
		memory[16'h3627] <= 8'ha2;
		memory[16'h3628] <= 8'h82;
		memory[16'h3629] <= 8'h18;
		memory[16'h362a] <= 8'hd4;
		memory[16'h362b] <= 8'hca;
		memory[16'h362c] <= 8'h53;
		memory[16'h362d] <= 8'h5;
		memory[16'h362e] <= 8'he3;
		memory[16'h362f] <= 8'h30;
		memory[16'h3630] <= 8'h14;
		memory[16'h3631] <= 8'hf3;
		memory[16'h3632] <= 8'hfd;
		memory[16'h3633] <= 8'h3b;
		memory[16'h3634] <= 8'h81;
		memory[16'h3635] <= 8'h83;
		memory[16'h3636] <= 8'h3b;
		memory[16'h3637] <= 8'ha5;
		memory[16'h3638] <= 8'h3f;
		memory[16'h3639] <= 8'h45;
		memory[16'h363a] <= 8'hd0;
		memory[16'h363b] <= 8'h9f;
		memory[16'h363c] <= 8'h4;
		memory[16'h363d] <= 8'h92;
		memory[16'h363e] <= 8'h8c;
		memory[16'h363f] <= 8'h56;
		memory[16'h3640] <= 8'h66;
		memory[16'h3641] <= 8'h9b;
		memory[16'h3642] <= 8'h49;
		memory[16'h3643] <= 8'h9b;
		memory[16'h3644] <= 8'hed;
		memory[16'h3645] <= 8'hc8;
		memory[16'h3646] <= 8'h3e;
		memory[16'h3647] <= 8'h6f;
		memory[16'h3648] <= 8'he1;
		memory[16'h3649] <= 8'h12;
		memory[16'h364a] <= 8'h39;
		memory[16'h364b] <= 8'h34;
		memory[16'h364c] <= 8'h17;
		memory[16'h364d] <= 8'h1d;
		memory[16'h364e] <= 8'h64;
		memory[16'h364f] <= 8'h2b;
		memory[16'h3650] <= 8'h10;
		memory[16'h3651] <= 8'h62;
		memory[16'h3652] <= 8'h66;
		memory[16'h3653] <= 8'h91;
		memory[16'h3654] <= 8'he5;
		memory[16'h3655] <= 8'ha1;
		memory[16'h3656] <= 8'h36;
		memory[16'h3657] <= 8'h24;
		memory[16'h3658] <= 8'he7;
		memory[16'h3659] <= 8'h7;
		memory[16'h365a] <= 8'hc3;
		memory[16'h365b] <= 8'heb;
		memory[16'h365c] <= 8'h99;
		memory[16'h365d] <= 8'h4f;
		memory[16'h365e] <= 8'h42;
		memory[16'h365f] <= 8'hff;
		memory[16'h3660] <= 8'hea;
		memory[16'h3661] <= 8'h8b;
		memory[16'h3662] <= 8'h9a;
		memory[16'h3663] <= 8'hd7;
		memory[16'h3664] <= 8'h54;
		memory[16'h3665] <= 8'hd8;
		memory[16'h3666] <= 8'h47;
		memory[16'h3667] <= 8'h35;
		memory[16'h3668] <= 8'heb;
		memory[16'h3669] <= 8'h80;
		memory[16'h366a] <= 8'h69;
		memory[16'h366b] <= 8'h2;
		memory[16'h366c] <= 8'h9d;
		memory[16'h366d] <= 8'hce;
		memory[16'h366e] <= 8'h2e;
		memory[16'h366f] <= 8'had;
		memory[16'h3670] <= 8'h30;
		memory[16'h3671] <= 8'h94;
		memory[16'h3672] <= 8'h3f;
		memory[16'h3673] <= 8'h15;
		memory[16'h3674] <= 8'h36;
		memory[16'h3675] <= 8'h75;
		memory[16'h3676] <= 8'h39;
		memory[16'h3677] <= 8'h1d;
		memory[16'h3678] <= 8'h7c;
		memory[16'h3679] <= 8'hfc;
		memory[16'h367a] <= 8'h8;
		memory[16'h367b] <= 8'h15;
		memory[16'h367c] <= 8'h4b;
		memory[16'h367d] <= 8'h4a;
		memory[16'h367e] <= 8'h14;
		memory[16'h367f] <= 8'h35;
		memory[16'h3680] <= 8'hd6;
		memory[16'h3681] <= 8'haf;
		memory[16'h3682] <= 8'hd;
		memory[16'h3683] <= 8'h2a;
		memory[16'h3684] <= 8'h87;
		memory[16'h3685] <= 8'h54;
		memory[16'h3686] <= 8'h5f;
		memory[16'h3687] <= 8'h72;
		memory[16'h3688] <= 8'hd4;
		memory[16'h3689] <= 8'hc8;
		memory[16'h368a] <= 8'h75;
		memory[16'h368b] <= 8'h72;
		memory[16'h368c] <= 8'h96;
		memory[16'h368d] <= 8'ha3;
		memory[16'h368e] <= 8'h1f;
		memory[16'h368f] <= 8'hc6;
		memory[16'h3690] <= 8'h37;
		memory[16'h3691] <= 8'h5e;
		memory[16'h3692] <= 8'hdb;
		memory[16'h3693] <= 8'h6d;
		memory[16'h3694] <= 8'hd4;
		memory[16'h3695] <= 8'h14;
		memory[16'h3696] <= 8'h8a;
		memory[16'h3697] <= 8'h50;
		memory[16'h3698] <= 8'h10;
		memory[16'h3699] <= 8'h93;
		memory[16'h369a] <= 8'h66;
		memory[16'h369b] <= 8'h5b;
		memory[16'h369c] <= 8'hdd;
		memory[16'h369d] <= 8'h7a;
		memory[16'h369e] <= 8'h91;
		memory[16'h369f] <= 8'hb3;
		memory[16'h36a0] <= 8'h29;
		memory[16'h36a1] <= 8'h9e;
		memory[16'h36a2] <= 8'hdd;
		memory[16'h36a3] <= 8'hb1;
		memory[16'h36a4] <= 8'hf2;
		memory[16'h36a5] <= 8'h3c;
		memory[16'h36a6] <= 8'h23;
		memory[16'h36a7] <= 8'hc6;
		memory[16'h36a8] <= 8'h5;
		memory[16'h36a9] <= 8'h98;
		memory[16'h36aa] <= 8'h38;
		memory[16'h36ab] <= 8'h9b;
		memory[16'h36ac] <= 8'h3b;
		memory[16'h36ad] <= 8'h58;
		memory[16'h36ae] <= 8'h62;
		memory[16'h36af] <= 8'h73;
		memory[16'h36b0] <= 8'hb6;
		memory[16'h36b1] <= 8'h3d;
		memory[16'h36b2] <= 8'he0;
		memory[16'h36b3] <= 8'h8a;
		memory[16'h36b4] <= 8'h52;
		memory[16'h36b5] <= 8'h6b;
		memory[16'h36b6] <= 8'hdb;
		memory[16'h36b7] <= 8'h62;
		memory[16'h36b8] <= 8'hfe;
		memory[16'h36b9] <= 8'h41;
		memory[16'h36ba] <= 8'hbe;
		memory[16'h36bb] <= 8'hdb;
		memory[16'h36bc] <= 8'hbb;
		memory[16'h36bd] <= 8'h4f;
		memory[16'h36be] <= 8'h8f;
		memory[16'h36bf] <= 8'he5;
		memory[16'h36c0] <= 8'hed;
		memory[16'h36c1] <= 8'h6c;
		memory[16'h36c2] <= 8'h96;
		memory[16'h36c3] <= 8'hdf;
		memory[16'h36c4] <= 8'ha9;
		memory[16'h36c5] <= 8'hb9;
		memory[16'h36c6] <= 8'ha5;
		memory[16'h36c7] <= 8'hae;
		memory[16'h36c8] <= 8'h52;
		memory[16'h36c9] <= 8'hde;
		memory[16'h36ca] <= 8'h49;
		memory[16'h36cb] <= 8'h8d;
		memory[16'h36cc] <= 8'h36;
		memory[16'h36cd] <= 8'hab;
		memory[16'h36ce] <= 8'h0;
		memory[16'h36cf] <= 8'hec;
		memory[16'h36d0] <= 8'he9;
		memory[16'h36d1] <= 8'he1;
		memory[16'h36d2] <= 8'h77;
		memory[16'h36d3] <= 8'h3b;
		memory[16'h36d4] <= 8'h4c;
		memory[16'h36d5] <= 8'h52;
		memory[16'h36d6] <= 8'h9d;
		memory[16'h36d7] <= 8'h4a;
		memory[16'h36d8] <= 8'h93;
		memory[16'h36d9] <= 8'h5b;
		memory[16'h36da] <= 8'h25;
		memory[16'h36db] <= 8'h4e;
		memory[16'h36dc] <= 8'haa;
		memory[16'h36dd] <= 8'hb4;
		memory[16'h36de] <= 8'h33;
		memory[16'h36df] <= 8'h97;
		memory[16'h36e0] <= 8'h21;
		memory[16'h36e1] <= 8'hc9;
		memory[16'h36e2] <= 8'h76;
		memory[16'h36e3] <= 8'hca;
		memory[16'h36e4] <= 8'h83;
		memory[16'h36e5] <= 8'h1c;
		memory[16'h36e6] <= 8'h78;
		memory[16'h36e7] <= 8'hd5;
		memory[16'h36e8] <= 8'hfa;
		memory[16'h36e9] <= 8'hc1;
		memory[16'h36ea] <= 8'h62;
		memory[16'h36eb] <= 8'h30;
		memory[16'h36ec] <= 8'h6d;
		memory[16'h36ed] <= 8'h63;
		memory[16'h36ee] <= 8'h1c;
		memory[16'h36ef] <= 8'h56;
		memory[16'h36f0] <= 8'h44;
		memory[16'h36f1] <= 8'h93;
		memory[16'h36f2] <= 8'h91;
		memory[16'h36f3] <= 8'h90;
		memory[16'h36f4] <= 8'he5;
		memory[16'h36f5] <= 8'h2e;
		memory[16'h36f6] <= 8'hda;
		memory[16'h36f7] <= 8'h78;
		memory[16'h36f8] <= 8'h8a;
		memory[16'h36f9] <= 8'hff;
		memory[16'h36fa] <= 8'hc7;
		memory[16'h36fb] <= 8'h34;
		memory[16'h36fc] <= 8'hb4;
		memory[16'h36fd] <= 8'hfa;
		memory[16'h36fe] <= 8'hcc;
		memory[16'h36ff] <= 8'hd5;
		memory[16'h3700] <= 8'hc4;
		memory[16'h3701] <= 8'h42;
		memory[16'h3702] <= 8'h9f;
		memory[16'h3703] <= 8'h47;
		memory[16'h3704] <= 8'h5e;
		memory[16'h3705] <= 8'h17;
		memory[16'h3706] <= 8'h1c;
		memory[16'h3707] <= 8'h58;
		memory[16'h3708] <= 8'hd8;
		memory[16'h3709] <= 8'h7e;
		memory[16'h370a] <= 8'h88;
		memory[16'h370b] <= 8'h45;
		memory[16'h370c] <= 8'he1;
		memory[16'h370d] <= 8'ha5;
		memory[16'h370e] <= 8'h9b;
		memory[16'h370f] <= 8'h25;
		memory[16'h3710] <= 8'h38;
		memory[16'h3711] <= 8'h2c;
		memory[16'h3712] <= 8'hb5;
		memory[16'h3713] <= 8'h1e;
		memory[16'h3714] <= 8'h5b;
		memory[16'h3715] <= 8'h8f;
		memory[16'h3716] <= 8'h96;
		memory[16'h3717] <= 8'he5;
		memory[16'h3718] <= 8'h8f;
		memory[16'h3719] <= 8'h5d;
		memory[16'h371a] <= 8'h19;
		memory[16'h371b] <= 8'h43;
		memory[16'h371c] <= 8'h58;
		memory[16'h371d] <= 8'he5;
		memory[16'h371e] <= 8'h18;
		memory[16'h371f] <= 8'h1c;
		memory[16'h3720] <= 8'h28;
		memory[16'h3721] <= 8'hb7;
		memory[16'h3722] <= 8'h63;
		memory[16'h3723] <= 8'h86;
		memory[16'h3724] <= 8'hce;
		memory[16'h3725] <= 8'h7f;
		memory[16'h3726] <= 8'hdf;
		memory[16'h3727] <= 8'ha6;
		memory[16'h3728] <= 8'hfd;
		memory[16'h3729] <= 8'h67;
		memory[16'h372a] <= 8'hec;
		memory[16'h372b] <= 8'hdf;
		memory[16'h372c] <= 8'hc;
		memory[16'h372d] <= 8'h87;
		memory[16'h372e] <= 8'h4;
		memory[16'h372f] <= 8'h45;
		memory[16'h3730] <= 8'hb4;
		memory[16'h3731] <= 8'hba;
		memory[16'h3732] <= 8'h63;
		memory[16'h3733] <= 8'hf;
		memory[16'h3734] <= 8'h49;
		memory[16'h3735] <= 8'hf9;
		memory[16'h3736] <= 8'hf4;
		memory[16'h3737] <= 8'hd8;
		memory[16'h3738] <= 8'h57;
		memory[16'h3739] <= 8'hd;
		memory[16'h373a] <= 8'h1b;
		memory[16'h373b] <= 8'haf;
		memory[16'h373c] <= 8'hf3;
		memory[16'h373d] <= 8'h33;
		memory[16'h373e] <= 8'hcb;
		memory[16'h373f] <= 8'h1b;
		memory[16'h3740] <= 8'hea;
		memory[16'h3741] <= 8'h2e;
		memory[16'h3742] <= 8'ha1;
		memory[16'h3743] <= 8'hb8;
		memory[16'h3744] <= 8'had;
		memory[16'h3745] <= 8'h80;
		memory[16'h3746] <= 8'h5f;
		memory[16'h3747] <= 8'haa;
		memory[16'h3748] <= 8'he8;
		memory[16'h3749] <= 8'h4b;
		memory[16'h374a] <= 8'h89;
		memory[16'h374b] <= 8'hf4;
		memory[16'h374c] <= 8'hd2;
		memory[16'h374d] <= 8'h8e;
		memory[16'h374e] <= 8'h39;
		memory[16'h374f] <= 8'h86;
		memory[16'h3750] <= 8'h48;
		memory[16'h3751] <= 8'h9c;
		memory[16'h3752] <= 8'h95;
		memory[16'h3753] <= 8'h91;
		memory[16'h3754] <= 8'h96;
		memory[16'h3755] <= 8'h89;
		memory[16'h3756] <= 8'h6a;
		memory[16'h3757] <= 8'hed;
		memory[16'h3758] <= 8'h97;
		memory[16'h3759] <= 8'h85;
		memory[16'h375a] <= 8'h9c;
		memory[16'h375b] <= 8'h8a;
		memory[16'h375c] <= 8'hb9;
		memory[16'h375d] <= 8'h67;
		memory[16'h375e] <= 8'ha5;
		memory[16'h375f] <= 8'ha3;
		memory[16'h3760] <= 8'h95;
		memory[16'h3761] <= 8'h46;
		memory[16'h3762] <= 8'h5c;
		memory[16'h3763] <= 8'h42;
		memory[16'h3764] <= 8'hc7;
		memory[16'h3765] <= 8'hbb;
		memory[16'h3766] <= 8'hec;
		memory[16'h3767] <= 8'haf;
		memory[16'h3768] <= 8'h6;
		memory[16'h3769] <= 8'h76;
		memory[16'h376a] <= 8'ha3;
		memory[16'h376b] <= 8'hd8;
		memory[16'h376c] <= 8'h4;
		memory[16'h376d] <= 8'hdd;
		memory[16'h376e] <= 8'h5f;
		memory[16'h376f] <= 8'h4c;
		memory[16'h3770] <= 8'h79;
		memory[16'h3771] <= 8'hf4;
		memory[16'h3772] <= 8'hdd;
		memory[16'h3773] <= 8'hf;
		memory[16'h3774] <= 8'h7e;
		memory[16'h3775] <= 8'h47;
		memory[16'h3776] <= 8'hfc;
		memory[16'h3777] <= 8'h15;
		memory[16'h3778] <= 8'hcd;
		memory[16'h3779] <= 8'h98;
		memory[16'h377a] <= 8'h9f;
		memory[16'h377b] <= 8'h86;
		memory[16'h377c] <= 8'hff;
		memory[16'h377d] <= 8'h44;
		memory[16'h377e] <= 8'h29;
		memory[16'h377f] <= 8'h94;
		memory[16'h3780] <= 8'h8a;
		memory[16'h3781] <= 8'h85;
		memory[16'h3782] <= 8'hd6;
		memory[16'h3783] <= 8'h51;
		memory[16'h3784] <= 8'h40;
		memory[16'h3785] <= 8'hc3;
		memory[16'h3786] <= 8'h0;
		memory[16'h3787] <= 8'h46;
		memory[16'h3788] <= 8'h39;
		memory[16'h3789] <= 8'ha4;
		memory[16'h378a] <= 8'h1f;
		memory[16'h378b] <= 8'h3d;
		memory[16'h378c] <= 8'h81;
		memory[16'h378d] <= 8'h7e;
		memory[16'h378e] <= 8'h89;
		memory[16'h378f] <= 8'hfa;
		memory[16'h3790] <= 8'h72;
		memory[16'h3791] <= 8'h66;
		memory[16'h3792] <= 8'ha;
		memory[16'h3793] <= 8'hf0;
		memory[16'h3794] <= 8'hae;
		memory[16'h3795] <= 8'h6;
		memory[16'h3796] <= 8'h5;
		memory[16'h3797] <= 8'h7b;
		memory[16'h3798] <= 8'h9f;
		memory[16'h3799] <= 8'ha4;
		memory[16'h379a] <= 8'h1;
		memory[16'h379b] <= 8'h9e;
		memory[16'h379c] <= 8'he8;
		memory[16'h379d] <= 8'h2a;
		memory[16'h379e] <= 8'h33;
		memory[16'h379f] <= 8'h73;
		memory[16'h37a0] <= 8'hb0;
		memory[16'h37a1] <= 8'h9;
		memory[16'h37a2] <= 8'hc4;
		memory[16'h37a3] <= 8'hf0;
		memory[16'h37a4] <= 8'hcc;
		memory[16'h37a5] <= 8'hc5;
		memory[16'h37a6] <= 8'h37;
		memory[16'h37a7] <= 8'h5;
		memory[16'h37a8] <= 8'h69;
		memory[16'h37a9] <= 8'h56;
		memory[16'h37aa] <= 8'h42;
		memory[16'h37ab] <= 8'hea;
		memory[16'h37ac] <= 8'hd4;
		memory[16'h37ad] <= 8'hcb;
		memory[16'h37ae] <= 8'he4;
		memory[16'h37af] <= 8'h46;
		memory[16'h37b0] <= 8'h32;
		memory[16'h37b1] <= 8'hee;
		memory[16'h37b2] <= 8'h37;
		memory[16'h37b3] <= 8'he0;
		memory[16'h37b4] <= 8'hf5;
		memory[16'h37b5] <= 8'h3c;
		memory[16'h37b6] <= 8'h5b;
		memory[16'h37b7] <= 8'h94;
		memory[16'h37b8] <= 8'he1;
		memory[16'h37b9] <= 8'h5c;
		memory[16'h37ba] <= 8'h32;
		memory[16'h37bb] <= 8'hc9;
		memory[16'h37bc] <= 8'h86;
		memory[16'h37bd] <= 8'h65;
		memory[16'h37be] <= 8'h3c;
		memory[16'h37bf] <= 8'h36;
		memory[16'h37c0] <= 8'h6f;
		memory[16'h37c1] <= 8'h1;
		memory[16'h37c2] <= 8'h27;
		memory[16'h37c3] <= 8'h3b;
		memory[16'h37c4] <= 8'hc6;
		memory[16'h37c5] <= 8'h5e;
		memory[16'h37c6] <= 8'h41;
		memory[16'h37c7] <= 8'h2f;
		memory[16'h37c8] <= 8'hb4;
		memory[16'h37c9] <= 8'h83;
		memory[16'h37ca] <= 8'h19;
		memory[16'h37cb] <= 8'h88;
		memory[16'h37cc] <= 8'h4f;
		memory[16'h37cd] <= 8'hfd;
		memory[16'h37ce] <= 8'hce;
		memory[16'h37cf] <= 8'h81;
		memory[16'h37d0] <= 8'hec;
		memory[16'h37d1] <= 8'h5;
		memory[16'h37d2] <= 8'h61;
		memory[16'h37d3] <= 8'he1;
		memory[16'h37d4] <= 8'h42;
		memory[16'h37d5] <= 8'hbc;
		memory[16'h37d6] <= 8'h75;
		memory[16'h37d7] <= 8'h23;
		memory[16'h37d8] <= 8'h18;
		memory[16'h37d9] <= 8'ha7;
		memory[16'h37da] <= 8'hec;
		memory[16'h37db] <= 8'h9e;
		memory[16'h37dc] <= 8'hd;
		memory[16'h37dd] <= 8'h29;
		memory[16'h37de] <= 8'hd5;
		memory[16'h37df] <= 8'h7c;
		memory[16'h37e0] <= 8'h2a;
		memory[16'h37e1] <= 8'hfc;
		memory[16'h37e2] <= 8'hb7;
		memory[16'h37e3] <= 8'hf0;
		memory[16'h37e4] <= 8'h5a;
		memory[16'h37e5] <= 8'hf8;
		memory[16'h37e6] <= 8'h1f;
		memory[16'h37e7] <= 8'he;
		memory[16'h37e8] <= 8'h7c;
		memory[16'h37e9] <= 8'h38;
		memory[16'h37ea] <= 8'h96;
		memory[16'h37eb] <= 8'hcb;
		memory[16'h37ec] <= 8'h35;
		memory[16'h37ed] <= 8'h64;
		memory[16'h37ee] <= 8'h4c;
		memory[16'h37ef] <= 8'h21;
		memory[16'h37f0] <= 8'h6a;
		memory[16'h37f1] <= 8'had;
		memory[16'h37f2] <= 8'h2;
		memory[16'h37f3] <= 8'hac;
		memory[16'h37f4] <= 8'h69;
		memory[16'h37f5] <= 8'h77;
		memory[16'h37f6] <= 8'hcf;
		memory[16'h37f7] <= 8'h81;
		memory[16'h37f8] <= 8'h1f;
		memory[16'h37f9] <= 8'hbb;
		memory[16'h37fa] <= 8'h1f;
		memory[16'h37fb] <= 8'h2c;
		memory[16'h37fc] <= 8'he4;
		memory[16'h37fd] <= 8'hf4;
		memory[16'h37fe] <= 8'ha8;
		memory[16'h37ff] <= 8'he;
		memory[16'h3800] <= 8'hf0;
		memory[16'h3801] <= 8'h5f;
		memory[16'h3802] <= 8'hfe;
		memory[16'h3803] <= 8'h4a;
		memory[16'h3804] <= 8'h58;
		memory[16'h3805] <= 8'h1d;
		memory[16'h3806] <= 8'h58;
		memory[16'h3807] <= 8'hd4;
		memory[16'h3808] <= 8'h55;
		memory[16'h3809] <= 8'hee;
		memory[16'h380a] <= 8'h9f;
		memory[16'h380b] <= 8'h8b;
		memory[16'h380c] <= 8'h53;
		memory[16'h380d] <= 8'heb;
		memory[16'h380e] <= 8'hac;
		memory[16'h380f] <= 8'hbd;
		memory[16'h3810] <= 8'h98;
		memory[16'h3811] <= 8'haf;
		memory[16'h3812] <= 8'h69;
		memory[16'h3813] <= 8'h1;
		memory[16'h3814] <= 8'h26;
		memory[16'h3815] <= 8'h38;
		memory[16'h3816] <= 8'h82;
		memory[16'h3817] <= 8'h45;
		memory[16'h3818] <= 8'hf3;
		memory[16'h3819] <= 8'ha1;
		memory[16'h381a] <= 8'h71;
		memory[16'h381b] <= 8'hd8;
		memory[16'h381c] <= 8'h96;
		memory[16'h381d] <= 8'h19;
		memory[16'h381e] <= 8'he6;
		memory[16'h381f] <= 8'h86;
		memory[16'h3820] <= 8'h79;
		memory[16'h3821] <= 8'he5;
		memory[16'h3822] <= 8'hd1;
		memory[16'h3823] <= 8'hd1;
		memory[16'h3824] <= 8'h2;
		memory[16'h3825] <= 8'h29;
		memory[16'h3826] <= 8'ha5;
		memory[16'h3827] <= 8'h58;
		memory[16'h3828] <= 8'h18;
		memory[16'h3829] <= 8'h44;
		memory[16'h382a] <= 8'he3;
		memory[16'h382b] <= 8'h6b;
		memory[16'h382c] <= 8'h2f;
		memory[16'h382d] <= 8'h8f;
		memory[16'h382e] <= 8'h28;
		memory[16'h382f] <= 8'hc7;
		memory[16'h3830] <= 8'h3e;
		memory[16'h3831] <= 8'h91;
		memory[16'h3832] <= 8'hc8;
		memory[16'h3833] <= 8'h65;
		memory[16'h3834] <= 8'hc9;
		memory[16'h3835] <= 8'h4a;
		memory[16'h3836] <= 8'haa;
		memory[16'h3837] <= 8'hbc;
		memory[16'h3838] <= 8'heb;
		memory[16'h3839] <= 8'h1c;
		memory[16'h383a] <= 8'h94;
		memory[16'h383b] <= 8'h81;
		memory[16'h383c] <= 8'h35;
		memory[16'h383d] <= 8'h7b;
		memory[16'h383e] <= 8'h8;
		memory[16'h383f] <= 8'hae;
		memory[16'h3840] <= 8'h60;
		memory[16'h3841] <= 8'hd9;
		memory[16'h3842] <= 8'h7f;
		memory[16'h3843] <= 8'h62;
		memory[16'h3844] <= 8'h2;
		memory[16'h3845] <= 8'h24;
		memory[16'h3846] <= 8'hba;
		memory[16'h3847] <= 8'h1a;
		memory[16'h3848] <= 8'h68;
		memory[16'h3849] <= 8'h9d;
		memory[16'h384a] <= 8'h85;
		memory[16'h384b] <= 8'h97;
		memory[16'h384c] <= 8'h2d;
		memory[16'h384d] <= 8'had;
		memory[16'h384e] <= 8'h5e;
		memory[16'h384f] <= 8'h6b;
		memory[16'h3850] <= 8'h3e;
		memory[16'h3851] <= 8'h26;
		memory[16'h3852] <= 8'hd0;
		memory[16'h3853] <= 8'h7;
		memory[16'h3854] <= 8'h70;
		memory[16'h3855] <= 8'h7b;
		memory[16'h3856] <= 8'hc4;
		memory[16'h3857] <= 8'h5c;
		memory[16'h3858] <= 8'h97;
		memory[16'h3859] <= 8'h58;
		memory[16'h385a] <= 8'hdd;
		memory[16'h385b] <= 8'hcc;
		memory[16'h385c] <= 8'hd3;
		memory[16'h385d] <= 8'he5;
		memory[16'h385e] <= 8'h7b;
		memory[16'h385f] <= 8'h33;
		memory[16'h3860] <= 8'hbe;
		memory[16'h3861] <= 8'hfa;
		memory[16'h3862] <= 8'h96;
		memory[16'h3863] <= 8'hc1;
		memory[16'h3864] <= 8'h1f;
		memory[16'h3865] <= 8'h50;
		memory[16'h3866] <= 8'hdb;
		memory[16'h3867] <= 8'h87;
		memory[16'h3868] <= 8'hee;
		memory[16'h3869] <= 8'h61;
		memory[16'h386a] <= 8'h1f;
		memory[16'h386b] <= 8'h1b;
		memory[16'h386c] <= 8'he;
		memory[16'h386d] <= 8'h7d;
		memory[16'h386e] <= 8'h86;
		memory[16'h386f] <= 8'h4d;
		memory[16'h3870] <= 8'ha4;
		memory[16'h3871] <= 8'h57;
		memory[16'h3872] <= 8'h54;
		memory[16'h3873] <= 8'h14;
		memory[16'h3874] <= 8'hd2;
		memory[16'h3875] <= 8'h18;
		memory[16'h3876] <= 8'h70;
		memory[16'h3877] <= 8'h69;
		memory[16'h3878] <= 8'h71;
		memory[16'h3879] <= 8'h4e;
		memory[16'h387a] <= 8'h35;
		memory[16'h387b] <= 8'h44;
		memory[16'h387c] <= 8'h33;
		memory[16'h387d] <= 8'hb0;
		memory[16'h387e] <= 8'h78;
		memory[16'h387f] <= 8'hf2;
		memory[16'h3880] <= 8'hab;
		memory[16'h3881] <= 8'he;
		memory[16'h3882] <= 8'hb3;
		memory[16'h3883] <= 8'hca;
		memory[16'h3884] <= 8'h5e;
		memory[16'h3885] <= 8'h8e;
		memory[16'h3886] <= 8'h51;
		memory[16'h3887] <= 8'h4c;
		memory[16'h3888] <= 8'hef;
		memory[16'h3889] <= 8'h70;
		memory[16'h388a] <= 8'h67;
		memory[16'h388b] <= 8'hfe;
		memory[16'h388c] <= 8'hee;
		memory[16'h388d] <= 8'hee;
		memory[16'h388e] <= 8'h4b;
		memory[16'h388f] <= 8'h92;
		memory[16'h3890] <= 8'h45;
		memory[16'h3891] <= 8'h9f;
		memory[16'h3892] <= 8'ha6;
		memory[16'h3893] <= 8'h17;
		memory[16'h3894] <= 8'hb8;
		memory[16'h3895] <= 8'h17;
		memory[16'h3896] <= 8'h80;
		memory[16'h3897] <= 8'h29;
		memory[16'h3898] <= 8'h65;
		memory[16'h3899] <= 8'hb5;
		memory[16'h389a] <= 8'h6d;
		memory[16'h389b] <= 8'h98;
		memory[16'h389c] <= 8'h66;
		memory[16'h389d] <= 8'he5;
		memory[16'h389e] <= 8'h8a;
		memory[16'h389f] <= 8'h11;
		memory[16'h38a0] <= 8'hf3;
		memory[16'h38a1] <= 8'h3d;
		memory[16'h38a2] <= 8'hdb;
		memory[16'h38a3] <= 8'h52;
		memory[16'h38a4] <= 8'hcc;
		memory[16'h38a5] <= 8'h2c;
		memory[16'h38a6] <= 8'h9e;
		memory[16'h38a7] <= 8'hbb;
		memory[16'h38a8] <= 8'h9d;
		memory[16'h38a9] <= 8'h6;
		memory[16'h38aa] <= 8'hb9;
		memory[16'h38ab] <= 8'h8b;
		memory[16'h38ac] <= 8'hf4;
		memory[16'h38ad] <= 8'h4;
		memory[16'h38ae] <= 8'h1d;
		memory[16'h38af] <= 8'h39;
		memory[16'h38b0] <= 8'ha4;
		memory[16'h38b1] <= 8'hc3;
		memory[16'h38b2] <= 8'h50;
		memory[16'h38b3] <= 8'h5c;
		memory[16'h38b4] <= 8'hda;
		memory[16'h38b5] <= 8'hd0;
		memory[16'h38b6] <= 8'h85;
		memory[16'h38b7] <= 8'h3f;
		memory[16'h38b8] <= 8'h85;
		memory[16'h38b9] <= 8'hf2;
		memory[16'h38ba] <= 8'hd8;
		memory[16'h38bb] <= 8'heb;
		memory[16'h38bc] <= 8'hd8;
		memory[16'h38bd] <= 8'h62;
		memory[16'h38be] <= 8'hfc;
		memory[16'h38bf] <= 8'hcb;
		memory[16'h38c0] <= 8'ha0;
		memory[16'h38c1] <= 8'hd7;
		memory[16'h38c2] <= 8'h1d;
		memory[16'h38c3] <= 8'h6c;
		memory[16'h38c4] <= 8'h4;
		memory[16'h38c5] <= 8'hbc;
		memory[16'h38c6] <= 8'h27;
		memory[16'h38c7] <= 8'ha1;
		memory[16'h38c8] <= 8'hc2;
		memory[16'h38c9] <= 8'he1;
		memory[16'h38ca] <= 8'h2c;
		memory[16'h38cb] <= 8'hb6;
		memory[16'h38cc] <= 8'he5;
		memory[16'h38cd] <= 8'h49;
		memory[16'h38ce] <= 8'hef;
		memory[16'h38cf] <= 8'h89;
		memory[16'h38d0] <= 8'hc;
		memory[16'h38d1] <= 8'h3f;
		memory[16'h38d2] <= 8'he5;
		memory[16'h38d3] <= 8'he7;
		memory[16'h38d4] <= 8'hf;
		memory[16'h38d5] <= 8'h6a;
		memory[16'h38d6] <= 8'h26;
		memory[16'h38d7] <= 8'h94;
		memory[16'h38d8] <= 8'h5d;
		memory[16'h38d9] <= 8'hfe;
		memory[16'h38da] <= 8'h80;
		memory[16'h38db] <= 8'h35;
		memory[16'h38dc] <= 8'h61;
		memory[16'h38dd] <= 8'h7c;
		memory[16'h38de] <= 8'h0;
		memory[16'h38df] <= 8'h1;
		memory[16'h38e0] <= 8'h54;
		memory[16'h38e1] <= 8'h1e;
		memory[16'h38e2] <= 8'h6d;
		memory[16'h38e3] <= 8'h58;
		memory[16'h38e4] <= 8'hda;
		memory[16'h38e5] <= 8'h94;
		memory[16'h38e6] <= 8'hf9;
		memory[16'h38e7] <= 8'h9c;
		memory[16'h38e8] <= 8'h75;
		memory[16'h38e9] <= 8'h25;
		memory[16'h38ea] <= 8'h52;
		memory[16'h38eb] <= 8'h5b;
		memory[16'h38ec] <= 8'h6e;
		memory[16'h38ed] <= 8'h41;
		memory[16'h38ee] <= 8'he4;
		memory[16'h38ef] <= 8'h7a;
		memory[16'h38f0] <= 8'h80;
		memory[16'h38f1] <= 8'hca;
		memory[16'h38f2] <= 8'h61;
		memory[16'h38f3] <= 8'h8f;
		memory[16'h38f4] <= 8'h34;
		memory[16'h38f5] <= 8'h88;
		memory[16'h38f6] <= 8'h23;
		memory[16'h38f7] <= 8'h91;
		memory[16'h38f8] <= 8'h86;
		memory[16'h38f9] <= 8'ha3;
		memory[16'h38fa] <= 8'hc6;
		memory[16'h38fb] <= 8'he7;
		memory[16'h38fc] <= 8'h20;
		memory[16'h38fd] <= 8'hc7;
		memory[16'h38fe] <= 8'he8;
		memory[16'h38ff] <= 8'h74;
		memory[16'h3900] <= 8'he5;
		memory[16'h3901] <= 8'h55;
		memory[16'h3902] <= 8'hcc;
		memory[16'h3903] <= 8'hbf;
		memory[16'h3904] <= 8'hea;
		memory[16'h3905] <= 8'hc5;
		memory[16'h3906] <= 8'h5b;
		memory[16'h3907] <= 8'h5f;
		memory[16'h3908] <= 8'hea;
		memory[16'h3909] <= 8'had;
		memory[16'h390a] <= 8'hba;
		memory[16'h390b] <= 8'h58;
		memory[16'h390c] <= 8'hee;
		memory[16'h390d] <= 8'h9f;
		memory[16'h390e] <= 8'hd2;
		memory[16'h390f] <= 8'h6e;
		memory[16'h3910] <= 8'h69;
		memory[16'h3911] <= 8'h34;
		memory[16'h3912] <= 8'hfd;
		memory[16'h3913] <= 8'h9d;
		memory[16'h3914] <= 8'hbc;
		memory[16'h3915] <= 8'h20;
		memory[16'h3916] <= 8'h2f;
		memory[16'h3917] <= 8'h42;
		memory[16'h3918] <= 8'hc4;
		memory[16'h3919] <= 8'hf5;
		memory[16'h391a] <= 8'h2a;
		memory[16'h391b] <= 8'he4;
		memory[16'h391c] <= 8'hbc;
		memory[16'h391d] <= 8'h12;
		memory[16'h391e] <= 8'h58;
		memory[16'h391f] <= 8'ha1;
		memory[16'h3920] <= 8'h68;
		memory[16'h3921] <= 8'h24;
		memory[16'h3922] <= 8'h60;
		memory[16'h3923] <= 8'h52;
		memory[16'h3924] <= 8'he9;
		memory[16'h3925] <= 8'hbb;
		memory[16'h3926] <= 8'hb1;
		memory[16'h3927] <= 8'hd3;
		memory[16'h3928] <= 8'h68;
		memory[16'h3929] <= 8'h6c;
		memory[16'h392a] <= 8'h2b;
		memory[16'h392b] <= 8'h56;
		memory[16'h392c] <= 8'hb;
		memory[16'h392d] <= 8'hfd;
		memory[16'h392e] <= 8'hc4;
		memory[16'h392f] <= 8'h74;
		memory[16'h3930] <= 8'h31;
		memory[16'h3931] <= 8'hc1;
		memory[16'h3932] <= 8'h11;
		memory[16'h3933] <= 8'hed;
		memory[16'h3934] <= 8'he2;
		memory[16'h3935] <= 8'h40;
		memory[16'h3936] <= 8'h30;
		memory[16'h3937] <= 8'ha6;
		memory[16'h3938] <= 8'h36;
		memory[16'h3939] <= 8'h5a;
		memory[16'h393a] <= 8'h8a;
		memory[16'h393b] <= 8'hf2;
		memory[16'h393c] <= 8'h6c;
		memory[16'h393d] <= 8'he2;
		memory[16'h393e] <= 8'h94;
		memory[16'h393f] <= 8'hd4;
		memory[16'h3940] <= 8'h6;
		memory[16'h3941] <= 8'hf4;
		memory[16'h3942] <= 8'h26;
		memory[16'h3943] <= 8'hef;
		memory[16'h3944] <= 8'hb0;
		memory[16'h3945] <= 8'hd8;
		memory[16'h3946] <= 8'hc2;
		memory[16'h3947] <= 8'h18;
		memory[16'h3948] <= 8'h44;
		memory[16'h3949] <= 8'hed;
		memory[16'h394a] <= 8'h6f;
		memory[16'h394b] <= 8'h4f;
		memory[16'h394c] <= 8'hea;
		memory[16'h394d] <= 8'h33;
		memory[16'h394e] <= 8'hc3;
		memory[16'h394f] <= 8'h1c;
		memory[16'h3950] <= 8'hf5;
		memory[16'h3951] <= 8'hd4;
		memory[16'h3952] <= 8'h9;
		memory[16'h3953] <= 8'hd7;
		memory[16'h3954] <= 8'h15;
		memory[16'h3955] <= 8'h39;
		memory[16'h3956] <= 8'h7d;
		memory[16'h3957] <= 8'h4b;
		memory[16'h3958] <= 8'h93;
		memory[16'h3959] <= 8'h7;
		memory[16'h395a] <= 8'h3d;
		memory[16'h395b] <= 8'h0;
		memory[16'h395c] <= 8'he9;
		memory[16'h395d] <= 8'hd1;
		memory[16'h395e] <= 8'hd4;
		memory[16'h395f] <= 8'hef;
		memory[16'h3960] <= 8'hc6;
		memory[16'h3961] <= 8'hfb;
		memory[16'h3962] <= 8'hde;
		memory[16'h3963] <= 8'h76;
		memory[16'h3964] <= 8'hd3;
		memory[16'h3965] <= 8'ha0;
		memory[16'h3966] <= 8'h8e;
		memory[16'h3967] <= 8'h17;
		memory[16'h3968] <= 8'h8d;
		memory[16'h3969] <= 8'hfd;
		memory[16'h396a] <= 8'h66;
		memory[16'h396b] <= 8'h77;
		memory[16'h396c] <= 8'h31;
		memory[16'h396d] <= 8'h29;
		memory[16'h396e] <= 8'h93;
		memory[16'h396f] <= 8'h26;
		memory[16'h3970] <= 8'hfd;
		memory[16'h3971] <= 8'h9d;
		memory[16'h3972] <= 8'hfd;
		memory[16'h3973] <= 8'h12;
		memory[16'h3974] <= 8'hd6;
		memory[16'h3975] <= 8'h7a;
		memory[16'h3976] <= 8'h5d;
		memory[16'h3977] <= 8'h6a;
		memory[16'h3978] <= 8'h81;
		memory[16'h3979] <= 8'h9b;
		memory[16'h397a] <= 8'h6a;
		memory[16'h397b] <= 8'h6a;
		memory[16'h397c] <= 8'h6c;
		memory[16'h397d] <= 8'h3e;
		memory[16'h397e] <= 8'h59;
		memory[16'h397f] <= 8'h32;
		memory[16'h3980] <= 8'h39;
		memory[16'h3981] <= 8'h37;
		memory[16'h3982] <= 8'ha8;
		memory[16'h3983] <= 8'hc;
		memory[16'h3984] <= 8'hd7;
		memory[16'h3985] <= 8'h37;
		memory[16'h3986] <= 8'h23;
		memory[16'h3987] <= 8'h64;
		memory[16'h3988] <= 8'h34;
		memory[16'h3989] <= 8'h89;
		memory[16'h398a] <= 8'hdb;
		memory[16'h398b] <= 8'h65;
		memory[16'h398c] <= 8'hb2;
		memory[16'h398d] <= 8'h6f;
		memory[16'h398e] <= 8'h8b;
		memory[16'h398f] <= 8'hb0;
		memory[16'h3990] <= 8'hc;
		memory[16'h3991] <= 8'h88;
		memory[16'h3992] <= 8'hc2;
		memory[16'h3993] <= 8'he2;
		memory[16'h3994] <= 8'h2;
		memory[16'h3995] <= 8'h20;
		memory[16'h3996] <= 8'h4c;
		memory[16'h3997] <= 8'h83;
		memory[16'h3998] <= 8'hbb;
		memory[16'h3999] <= 8'hb6;
		memory[16'h399a] <= 8'hed;
		memory[16'h399b] <= 8'h27;
		memory[16'h399c] <= 8'hf5;
		memory[16'h399d] <= 8'h46;
		memory[16'h399e] <= 8'h5a;
		memory[16'h399f] <= 8'h2e;
		memory[16'h39a0] <= 8'h7d;
		memory[16'h39a1] <= 8'h2;
		memory[16'h39a2] <= 8'h3b;
		memory[16'h39a3] <= 8'h54;
		memory[16'h39a4] <= 8'h39;
		memory[16'h39a5] <= 8'h5e;
		memory[16'h39a6] <= 8'hb8;
		memory[16'h39a7] <= 8'h6e;
		memory[16'h39a8] <= 8'he8;
		memory[16'h39a9] <= 8'h94;
		memory[16'h39aa] <= 8'hd3;
		memory[16'h39ab] <= 8'h9a;
		memory[16'h39ac] <= 8'h3;
		memory[16'h39ad] <= 8'h5f;
		memory[16'h39ae] <= 8'h4a;
		memory[16'h39af] <= 8'hf;
		memory[16'h39b0] <= 8'he7;
		memory[16'h39b1] <= 8'hd;
		memory[16'h39b2] <= 8'hf1;
		memory[16'h39b3] <= 8'hea;
		memory[16'h39b4] <= 8'h2d;
		memory[16'h39b5] <= 8'h3e;
		memory[16'h39b6] <= 8'h6d;
		memory[16'h39b7] <= 8'he8;
		memory[16'h39b8] <= 8'hf4;
		memory[16'h39b9] <= 8'h5b;
		memory[16'h39ba] <= 8'hf;
		memory[16'h39bb] <= 8'he9;
		memory[16'h39bc] <= 8'ha1;
		memory[16'h39bd] <= 8'h69;
		memory[16'h39be] <= 8'h18;
		memory[16'h39bf] <= 8'h1f;
		memory[16'h39c0] <= 8'h6c;
		memory[16'h39c1] <= 8'h53;
		memory[16'h39c2] <= 8'h73;
		memory[16'h39c3] <= 8'ha5;
		memory[16'h39c4] <= 8'hb1;
		memory[16'h39c5] <= 8'h2c;
		memory[16'h39c6] <= 8'h13;
		memory[16'h39c7] <= 8'h99;
		memory[16'h39c8] <= 8'hc0;
		memory[16'h39c9] <= 8'he7;
		memory[16'h39ca] <= 8'h34;
		memory[16'h39cb] <= 8'hc3;
		memory[16'h39cc] <= 8'h46;
		memory[16'h39cd] <= 8'h7e;
		memory[16'h39ce] <= 8'hd2;
		memory[16'h39cf] <= 8'h2d;
		memory[16'h39d0] <= 8'h8b;
		memory[16'h39d1] <= 8'hc3;
		memory[16'h39d2] <= 8'h17;
		memory[16'h39d3] <= 8'hb8;
		memory[16'h39d4] <= 8'h1;
		memory[16'h39d5] <= 8'h85;
		memory[16'h39d6] <= 8'ha0;
		memory[16'h39d7] <= 8'hf6;
		memory[16'h39d8] <= 8'he0;
		memory[16'h39d9] <= 8'hb0;
		memory[16'h39da] <= 8'hdf;
		memory[16'h39db] <= 8'h81;
		memory[16'h39dc] <= 8'h19;
		memory[16'h39dd] <= 8'hf7;
		memory[16'h39de] <= 8'ha0;
		memory[16'h39df] <= 8'h85;
		memory[16'h39e0] <= 8'h4a;
		memory[16'h39e1] <= 8'h14;
		memory[16'h39e2] <= 8'h2b;
		memory[16'h39e3] <= 8'hfc;
		memory[16'h39e4] <= 8'h40;
		memory[16'h39e5] <= 8'h3e;
		memory[16'h39e6] <= 8'h95;
		memory[16'h39e7] <= 8'h0;
		memory[16'h39e8] <= 8'h25;
		memory[16'h39e9] <= 8'hc9;
		memory[16'h39ea] <= 8'hc3;
		memory[16'h39eb] <= 8'h6b;
		memory[16'h39ec] <= 8'h48;
		memory[16'h39ed] <= 8'h95;
		memory[16'h39ee] <= 8'h99;
		memory[16'h39ef] <= 8'hd3;
		memory[16'h39f0] <= 8'h58;
		memory[16'h39f1] <= 8'hb0;
		memory[16'h39f2] <= 8'h8c;
		memory[16'h39f3] <= 8'h5a;
		memory[16'h39f4] <= 8'h35;
		memory[16'h39f5] <= 8'h2c;
		memory[16'h39f6] <= 8'h50;
		memory[16'h39f7] <= 8'h15;
		memory[16'h39f8] <= 8'hdc;
		memory[16'h39f9] <= 8'h2f;
		memory[16'h39fa] <= 8'h97;
		memory[16'h39fb] <= 8'hf6;
		memory[16'h39fc] <= 8'h27;
		memory[16'h39fd] <= 8'h37;
		memory[16'h39fe] <= 8'h7b;
		memory[16'h39ff] <= 8'h71;
		memory[16'h3a00] <= 8'h4b;
		memory[16'h3a01] <= 8'ha6;
		memory[16'h3a02] <= 8'h6d;
		memory[16'h3a03] <= 8'h8b;
		memory[16'h3a04] <= 8'he5;
		memory[16'h3a05] <= 8'h3;
		memory[16'h3a06] <= 8'h8b;
		memory[16'h3a07] <= 8'ha;
		memory[16'h3a08] <= 8'hcc;
		memory[16'h3a09] <= 8'h4e;
		memory[16'h3a0a] <= 8'h76;
		memory[16'h3a0b] <= 8'h14;
		memory[16'h3a0c] <= 8'he3;
		memory[16'h3a0d] <= 8'hf;
		memory[16'h3a0e] <= 8'he8;
		memory[16'h3a0f] <= 8'h3c;
		memory[16'h3a10] <= 8'hbf;
		memory[16'h3a11] <= 8'h74;
		memory[16'h3a12] <= 8'h96;
		memory[16'h3a13] <= 8'hf5;
		memory[16'h3a14] <= 8'ha0;
		memory[16'h3a15] <= 8'he6;
		memory[16'h3a16] <= 8'ha;
		memory[16'h3a17] <= 8'h7d;
		memory[16'h3a18] <= 8'h15;
		memory[16'h3a19] <= 8'ha1;
		memory[16'h3a1a] <= 8'h73;
		memory[16'h3a1b] <= 8'h3c;
		memory[16'h3a1c] <= 8'hd9;
		memory[16'h3a1d] <= 8'hee;
		memory[16'h3a1e] <= 8'hae;
		memory[16'h3a1f] <= 8'h24;
		memory[16'h3a20] <= 8'h95;
		memory[16'h3a21] <= 8'h1b;
		memory[16'h3a22] <= 8'hb0;
		memory[16'h3a23] <= 8'h7a;
		memory[16'h3a24] <= 8'h1e;
		memory[16'h3a25] <= 8'h3b;
		memory[16'h3a26] <= 8'h84;
		memory[16'h3a27] <= 8'heb;
		memory[16'h3a28] <= 8'h8a;
		memory[16'h3a29] <= 8'hfa;
		memory[16'h3a2a] <= 8'hff;
		memory[16'h3a2b] <= 8'h6d;
		memory[16'h3a2c] <= 8'h9;
		memory[16'h3a2d] <= 8'he7;
		memory[16'h3a2e] <= 8'ha9;
		memory[16'h3a2f] <= 8'hc9;
		memory[16'h3a30] <= 8'h5b;
		memory[16'h3a31] <= 8'h3f;
		memory[16'h3a32] <= 8'hbe;
		memory[16'h3a33] <= 8'hfc;
		memory[16'h3a34] <= 8'h25;
		memory[16'h3a35] <= 8'hc8;
		memory[16'h3a36] <= 8'h79;
		memory[16'h3a37] <= 8'h3b;
		memory[16'h3a38] <= 8'h6a;
		memory[16'h3a39] <= 8'hec;
		memory[16'h3a3a] <= 8'h77;
		memory[16'h3a3b] <= 8'h43;
		memory[16'h3a3c] <= 8'hda;
		memory[16'h3a3d] <= 8'h25;
		memory[16'h3a3e] <= 8'h67;
		memory[16'h3a3f] <= 8'h6f;
		memory[16'h3a40] <= 8'h41;
		memory[16'h3a41] <= 8'h17;
		memory[16'h3a42] <= 8'he9;
		memory[16'h3a43] <= 8'h5f;
		memory[16'h3a44] <= 8'h53;
		memory[16'h3a45] <= 8'h6e;
		memory[16'h3a46] <= 8'h4a;
		memory[16'h3a47] <= 8'hdd;
		memory[16'h3a48] <= 8'h68;
		memory[16'h3a49] <= 8'h4a;
		memory[16'h3a4a] <= 8'h4a;
		memory[16'h3a4b] <= 8'h72;
		memory[16'h3a4c] <= 8'h31;
		memory[16'h3a4d] <= 8'hf4;
		memory[16'h3a4e] <= 8'h3b;
		memory[16'h3a4f] <= 8'h8d;
		memory[16'h3a50] <= 8'h33;
		memory[16'h3a51] <= 8'hf9;
		memory[16'h3a52] <= 8'h89;
		memory[16'h3a53] <= 8'h59;
		memory[16'h3a54] <= 8'hc1;
		memory[16'h3a55] <= 8'h2;
		memory[16'h3a56] <= 8'h94;
		memory[16'h3a57] <= 8'h2b;
		memory[16'h3a58] <= 8'hee;
		memory[16'h3a59] <= 8'hb;
		memory[16'h3a5a] <= 8'h6e;
		memory[16'h3a5b] <= 8'hc8;
		memory[16'h3a5c] <= 8'h31;
		memory[16'h3a5d] <= 8'hd6;
		memory[16'h3a5e] <= 8'h38;
		memory[16'h3a5f] <= 8'h72;
		memory[16'h3a60] <= 8'hed;
		memory[16'h3a61] <= 8'h21;
		memory[16'h3a62] <= 8'hd1;
		memory[16'h3a63] <= 8'h40;
		memory[16'h3a64] <= 8'h8f;
		memory[16'h3a65] <= 8'h1c;
		memory[16'h3a66] <= 8'h1d;
		memory[16'h3a67] <= 8'hf8;
		memory[16'h3a68] <= 8'h66;
		memory[16'h3a69] <= 8'h68;
		memory[16'h3a6a] <= 8'h6a;
		memory[16'h3a6b] <= 8'h97;
		memory[16'h3a6c] <= 8'h5c;
		memory[16'h3a6d] <= 8'ha5;
		memory[16'h3a6e] <= 8'h24;
		memory[16'h3a6f] <= 8'h8f;
		memory[16'h3a70] <= 8'h9e;
		memory[16'h3a71] <= 8'had;
		memory[16'h3a72] <= 8'he8;
		memory[16'h3a73] <= 8'h5f;
		memory[16'h3a74] <= 8'haf;
		memory[16'h3a75] <= 8'h7c;
		memory[16'h3a76] <= 8'h8b;
		memory[16'h3a77] <= 8'h9d;
		memory[16'h3a78] <= 8'h88;
		memory[16'h3a79] <= 8'hf9;
		memory[16'h3a7a] <= 8'h66;
		memory[16'h3a7b] <= 8'hb9;
		memory[16'h3a7c] <= 8'hcf;
		memory[16'h3a7d] <= 8'h9e;
		memory[16'h3a7e] <= 8'h2b;
		memory[16'h3a7f] <= 8'hbd;
		memory[16'h3a80] <= 8'hbf;
		memory[16'h3a81] <= 8'hfc;
		memory[16'h3a82] <= 8'hfd;
		memory[16'h3a83] <= 8'h4f;
		memory[16'h3a84] <= 8'h18;
		memory[16'h3a85] <= 8'h1b;
		memory[16'h3a86] <= 8'h47;
		memory[16'h3a87] <= 8'h7e;
		memory[16'h3a88] <= 8'h83;
		memory[16'h3a89] <= 8'hb1;
		memory[16'h3a8a] <= 8'h16;
		memory[16'h3a8b] <= 8'hdf;
		memory[16'h3a8c] <= 8'h56;
		memory[16'h3a8d] <= 8'h3a;
		memory[16'h3a8e] <= 8'h6e;
		memory[16'h3a8f] <= 8'hf4;
		memory[16'h3a90] <= 8'he8;
		memory[16'h3a91] <= 8'h57;
		memory[16'h3a92] <= 8'h53;
		memory[16'h3a93] <= 8'h97;
		memory[16'h3a94] <= 8'hd3;
		memory[16'h3a95] <= 8'hde;
		memory[16'h3a96] <= 8'h35;
		memory[16'h3a97] <= 8'h5b;
		memory[16'h3a98] <= 8'hd8;
		memory[16'h3a99] <= 8'h9b;
		memory[16'h3a9a] <= 8'h14;
		memory[16'h3a9b] <= 8'ha7;
		memory[16'h3a9c] <= 8'h39;
		memory[16'h3a9d] <= 8'h3f;
		memory[16'h3a9e] <= 8'h64;
		memory[16'h3a9f] <= 8'hf8;
		memory[16'h3aa0] <= 8'h3c;
		memory[16'h3aa1] <= 8'h62;
		memory[16'h3aa2] <= 8'h47;
		memory[16'h3aa3] <= 8'h54;
		memory[16'h3aa4] <= 8'h7d;
		memory[16'h3aa5] <= 8'h8e;
		memory[16'h3aa6] <= 8'hd3;
		memory[16'h3aa7] <= 8'h0;
		memory[16'h3aa8] <= 8'h3f;
		memory[16'h3aa9] <= 8'he9;
		memory[16'h3aaa] <= 8'hdf;
		memory[16'h3aab] <= 8'h95;
		memory[16'h3aac] <= 8'h23;
		memory[16'h3aad] <= 8'h4d;
		memory[16'h3aae] <= 8'h89;
		memory[16'h3aaf] <= 8'hb;
		memory[16'h3ab0] <= 8'ha4;
		memory[16'h3ab1] <= 8'hdd;
		memory[16'h3ab2] <= 8'ha3;
		memory[16'h3ab3] <= 8'h78;
		memory[16'h3ab4] <= 8'hbb;
		memory[16'h3ab5] <= 8'hd8;
		memory[16'h3ab6] <= 8'hd3;
		memory[16'h3ab7] <= 8'h93;
		memory[16'h3ab8] <= 8'h73;
		memory[16'h3ab9] <= 8'he8;
		memory[16'h3aba] <= 8'h3b;
		memory[16'h3abb] <= 8'hac;
		memory[16'h3abc] <= 8'h27;
		memory[16'h3abd] <= 8'h9f;
		memory[16'h3abe] <= 8'ha4;
		memory[16'h3abf] <= 8'h63;
		memory[16'h3ac0] <= 8'h1;
		memory[16'h3ac1] <= 8'hec;
		memory[16'h3ac2] <= 8'hb8;
		memory[16'h3ac3] <= 8'h7e;
		memory[16'h3ac4] <= 8'h7a;
		memory[16'h3ac5] <= 8'h8b;
		memory[16'h3ac6] <= 8'h7e;
		memory[16'h3ac7] <= 8'hba;
		memory[16'h3ac8] <= 8'h74;
		memory[16'h3ac9] <= 8'h5d;
		memory[16'h3aca] <= 8'h4f;
		memory[16'h3acb] <= 8'h97;
		memory[16'h3acc] <= 8'hab;
		memory[16'h3acd] <= 8'hd9;
		memory[16'h3ace] <= 8'ha3;
		memory[16'h3acf] <= 8'h4f;
		memory[16'h3ad0] <= 8'hb6;
		memory[16'h3ad1] <= 8'h46;
		memory[16'h3ad2] <= 8'hc7;
		memory[16'h3ad3] <= 8'h71;
		memory[16'h3ad4] <= 8'h1e;
		memory[16'h3ad5] <= 8'h9b;
		memory[16'h3ad6] <= 8'h5;
		memory[16'h3ad7] <= 8'h91;
		memory[16'h3ad8] <= 8'h83;
		memory[16'h3ad9] <= 8'h40;
		memory[16'h3ada] <= 8'h3d;
		memory[16'h3adb] <= 8'haa;
		memory[16'h3adc] <= 8'hdf;
		memory[16'h3add] <= 8'he1;
		memory[16'h3ade] <= 8'he;
		memory[16'h3adf] <= 8'he1;
		memory[16'h3ae0] <= 8'hcd;
		memory[16'h3ae1] <= 8'hc6;
		memory[16'h3ae2] <= 8'h5f;
		memory[16'h3ae3] <= 8'h48;
		memory[16'h3ae4] <= 8'h51;
		memory[16'h3ae5] <= 8'hde;
		memory[16'h3ae6] <= 8'h2;
		memory[16'h3ae7] <= 8'hc5;
		memory[16'h3ae8] <= 8'h3b;
		memory[16'h3ae9] <= 8'h51;
		memory[16'h3aea] <= 8'h5c;
		memory[16'h3aeb] <= 8'he6;
		memory[16'h3aec] <= 8'h2a;
		memory[16'h3aed] <= 8'hff;
		memory[16'h3aee] <= 8'h36;
		memory[16'h3aef] <= 8'he0;
		memory[16'h3af0] <= 8'h45;
		memory[16'h3af1] <= 8'hfd;
		memory[16'h3af2] <= 8'h52;
		memory[16'h3af3] <= 8'h63;
		memory[16'h3af4] <= 8'h98;
		memory[16'h3af5] <= 8'h57;
		memory[16'h3af6] <= 8'hf4;
		memory[16'h3af7] <= 8'h1b;
		memory[16'h3af8] <= 8'h97;
		memory[16'h3af9] <= 8'h31;
		memory[16'h3afa] <= 8'hc6;
		memory[16'h3afb] <= 8'h76;
		memory[16'h3afc] <= 8'h13;
		memory[16'h3afd] <= 8'hd4;
		memory[16'h3afe] <= 8'h57;
		memory[16'h3aff] <= 8'he0;
		memory[16'h3b00] <= 8'h9a;
		memory[16'h3b01] <= 8'hb7;
		memory[16'h3b02] <= 8'h28;
		memory[16'h3b03] <= 8'heb;
		memory[16'h3b04] <= 8'h95;
		memory[16'h3b05] <= 8'h2a;
		memory[16'h3b06] <= 8'hb0;
		memory[16'h3b07] <= 8'hd0;
		memory[16'h3b08] <= 8'h7c;
		memory[16'h3b09] <= 8'hc;
		memory[16'h3b0a] <= 8'hb7;
		memory[16'h3b0b] <= 8'ha6;
		memory[16'h3b0c] <= 8'hc;
		memory[16'h3b0d] <= 8'hed;
		memory[16'h3b0e] <= 8'h87;
		memory[16'h3b0f] <= 8'h51;
		memory[16'h3b10] <= 8'hea;
		memory[16'h3b11] <= 8'hd9;
		memory[16'h3b12] <= 8'hb5;
		memory[16'h3b13] <= 8'h83;
		memory[16'h3b14] <= 8'h30;
		memory[16'h3b15] <= 8'ha9;
		memory[16'h3b16] <= 8'h9e;
		memory[16'h3b17] <= 8'hc7;
		memory[16'h3b18] <= 8'hdb;
		memory[16'h3b19] <= 8'h64;
		memory[16'h3b1a] <= 8'h3d;
		memory[16'h3b1b] <= 8'hee;
		memory[16'h3b1c] <= 8'h38;
		memory[16'h3b1d] <= 8'h95;
		memory[16'h3b1e] <= 8'hce;
		memory[16'h3b1f] <= 8'hd2;
		memory[16'h3b20] <= 8'h4c;
		memory[16'h3b21] <= 8'hf7;
		memory[16'h3b22] <= 8'hbd;
		memory[16'h3b23] <= 8'he1;
		memory[16'h3b24] <= 8'h21;
		memory[16'h3b25] <= 8'h6d;
		memory[16'h3b26] <= 8'hb1;
		memory[16'h3b27] <= 8'h9d;
		memory[16'h3b28] <= 8'h7a;
		memory[16'h3b29] <= 8'h68;
		memory[16'h3b2a] <= 8'h44;
		memory[16'h3b2b] <= 8'h86;
		memory[16'h3b2c] <= 8'h55;
		memory[16'h3b2d] <= 8'hcb;
		memory[16'h3b2e] <= 8'hd7;
		memory[16'h3b2f] <= 8'h40;
		memory[16'h3b30] <= 8'ha4;
		memory[16'h3b31] <= 8'h8c;
		memory[16'h3b32] <= 8'hc3;
		memory[16'h3b33] <= 8'hd4;
		memory[16'h3b34] <= 8'h36;
		memory[16'h3b35] <= 8'h61;
		memory[16'h3b36] <= 8'h9b;
		memory[16'h3b37] <= 8'h11;
		memory[16'h3b38] <= 8'hc6;
		memory[16'h3b39] <= 8'hd8;
		memory[16'h3b3a] <= 8'hff;
		memory[16'h3b3b] <= 8'hfe;
		memory[16'h3b3c] <= 8'h6d;
		memory[16'h3b3d] <= 8'hcd;
		memory[16'h3b3e] <= 8'hd1;
		memory[16'h3b3f] <= 8'hb9;
		memory[16'h3b40] <= 8'hc4;
		memory[16'h3b41] <= 8'h8e;
		memory[16'h3b42] <= 8'h9a;
		memory[16'h3b43] <= 8'he6;
		memory[16'h3b44] <= 8'hfc;
		memory[16'h3b45] <= 8'h4c;
		memory[16'h3b46] <= 8'h83;
		memory[16'h3b47] <= 8'h76;
		memory[16'h3b48] <= 8'hb4;
		memory[16'h3b49] <= 8'hc7;
		memory[16'h3b4a] <= 8'hfc;
		memory[16'h3b4b] <= 8'ha;
		memory[16'h3b4c] <= 8'h92;
		memory[16'h3b4d] <= 8'hd3;
		memory[16'h3b4e] <= 8'h4a;
		memory[16'h3b4f] <= 8'h36;
		memory[16'h3b50] <= 8'h60;
		memory[16'h3b51] <= 8'hd;
		memory[16'h3b52] <= 8'ha;
		memory[16'h3b53] <= 8'h96;
		memory[16'h3b54] <= 8'h6e;
		memory[16'h3b55] <= 8'ha5;
		memory[16'h3b56] <= 8'ha7;
		memory[16'h3b57] <= 8'h34;
		memory[16'h3b58] <= 8'h7e;
		memory[16'h3b59] <= 8'ha6;
		memory[16'h3b5a] <= 8'h33;
		memory[16'h3b5b] <= 8'heb;
		memory[16'h3b5c] <= 8'h73;
		memory[16'h3b5d] <= 8'h4;
		memory[16'h3b5e] <= 8'ha5;
		memory[16'h3b5f] <= 8'h38;
		memory[16'h3b60] <= 8'h92;
		memory[16'h3b61] <= 8'h3f;
		memory[16'h3b62] <= 8'h1e;
		memory[16'h3b63] <= 8'h8e;
		memory[16'h3b64] <= 8'h8b;
		memory[16'h3b65] <= 8'ha1;
		memory[16'h3b66] <= 8'h4;
		memory[16'h3b67] <= 8'h40;
		memory[16'h3b68] <= 8'h69;
		memory[16'h3b69] <= 8'h0;
		memory[16'h3b6a] <= 8'h4a;
		memory[16'h3b6b] <= 8'hfb;
		memory[16'h3b6c] <= 8'hd4;
		memory[16'h3b6d] <= 8'h94;
		memory[16'h3b6e] <= 8'h32;
		memory[16'h3b6f] <= 8'h34;
		memory[16'h3b70] <= 8'ha1;
		memory[16'h3b71] <= 8'h3c;
		memory[16'h3b72] <= 8'hca;
		memory[16'h3b73] <= 8'hf;
		memory[16'h3b74] <= 8'he2;
		memory[16'h3b75] <= 8'h71;
		memory[16'h3b76] <= 8'h44;
		memory[16'h3b77] <= 8'h60;
		memory[16'h3b78] <= 8'h17;
		memory[16'h3b79] <= 8'h77;
		memory[16'h3b7a] <= 8'h4b;
		memory[16'h3b7b] <= 8'h8a;
		memory[16'h3b7c] <= 8'h7b;
		memory[16'h3b7d] <= 8'hf0;
		memory[16'h3b7e] <= 8'hc2;
		memory[16'h3b7f] <= 8'hd;
		memory[16'h3b80] <= 8'h30;
		memory[16'h3b81] <= 8'he0;
		memory[16'h3b82] <= 8'h9c;
		memory[16'h3b83] <= 8'hbb;
		memory[16'h3b84] <= 8'h82;
		memory[16'h3b85] <= 8'ha0;
		memory[16'h3b86] <= 8'hfb;
		memory[16'h3b87] <= 8'heb;
		memory[16'h3b88] <= 8'ha1;
		memory[16'h3b89] <= 8'h45;
		memory[16'h3b8a] <= 8'he6;
		memory[16'h3b8b] <= 8'h75;
		memory[16'h3b8c] <= 8'hd9;
		memory[16'h3b8d] <= 8'h18;
		memory[16'h3b8e] <= 8'ha9;
		memory[16'h3b8f] <= 8'h7a;
		memory[16'h3b90] <= 8'h55;
		memory[16'h3b91] <= 8'h73;
		memory[16'h3b92] <= 8'h8a;
		memory[16'h3b93] <= 8'h37;
		memory[16'h3b94] <= 8'he4;
		memory[16'h3b95] <= 8'hce;
		memory[16'h3b96] <= 8'h97;
		memory[16'h3b97] <= 8'hfb;
		memory[16'h3b98] <= 8'h45;
		memory[16'h3b99] <= 8'he2;
		memory[16'h3b9a] <= 8'h85;
		memory[16'h3b9b] <= 8'hc0;
		memory[16'h3b9c] <= 8'hd3;
		memory[16'h3b9d] <= 8'h48;
		memory[16'h3b9e] <= 8'hcd;
		memory[16'h3b9f] <= 8'h3;
		memory[16'h3ba0] <= 8'h28;
		memory[16'h3ba1] <= 8'h69;
		memory[16'h3ba2] <= 8'hbe;
		memory[16'h3ba3] <= 8'haa;
		memory[16'h3ba4] <= 8'ha;
		memory[16'h3ba5] <= 8'hba;
		memory[16'h3ba6] <= 8'h95;
		memory[16'h3ba7] <= 8'hab;
		memory[16'h3ba8] <= 8'hff;
		memory[16'h3ba9] <= 8'h7c;
		memory[16'h3baa] <= 8'h20;
		memory[16'h3bab] <= 8'hd9;
		memory[16'h3bac] <= 8'h94;
		memory[16'h3bad] <= 8'hc9;
		memory[16'h3bae] <= 8'h53;
		memory[16'h3baf] <= 8'he9;
		memory[16'h3bb0] <= 8'h3c;
		memory[16'h3bb1] <= 8'hdd;
		memory[16'h3bb2] <= 8'h20;
		memory[16'h3bb3] <= 8'h20;
		memory[16'h3bb4] <= 8'hab;
		memory[16'h3bb5] <= 8'hb7;
		memory[16'h3bb6] <= 8'h1b;
		memory[16'h3bb7] <= 8'hf0;
		memory[16'h3bb8] <= 8'h9a;
		memory[16'h3bb9] <= 8'ha0;
		memory[16'h3bba] <= 8'hb0;
		memory[16'h3bbb] <= 8'h6d;
		memory[16'h3bbc] <= 8'he8;
		memory[16'h3bbd] <= 8'h7e;
		memory[16'h3bbe] <= 8'h70;
		memory[16'h3bbf] <= 8'h11;
		memory[16'h3bc0] <= 8'he7;
		memory[16'h3bc1] <= 8'h2e;
		memory[16'h3bc2] <= 8'hbb;
		memory[16'h3bc3] <= 8'hf1;
		memory[16'h3bc4] <= 8'he8;
		memory[16'h3bc5] <= 8'h51;
		memory[16'h3bc6] <= 8'h9c;
		memory[16'h3bc7] <= 8'he8;
		memory[16'h3bc8] <= 8'hcd;
		memory[16'h3bc9] <= 8'hbc;
		memory[16'h3bca] <= 8'hc1;
		memory[16'h3bcb] <= 8'h61;
		memory[16'h3bcc] <= 8'h85;
		memory[16'h3bcd] <= 8'h14;
		memory[16'h3bce] <= 8'h4b;
		memory[16'h3bcf] <= 8'hc1;
		memory[16'h3bd0] <= 8'hf2;
		memory[16'h3bd1] <= 8'h6b;
		memory[16'h3bd2] <= 8'he1;
		memory[16'h3bd3] <= 8'h9d;
		memory[16'h3bd4] <= 8'h23;
		memory[16'h3bd5] <= 8'hfc;
		memory[16'h3bd6] <= 8'h8e;
		memory[16'h3bd7] <= 8'hbd;
		memory[16'h3bd8] <= 8'h9d;
		memory[16'h3bd9] <= 8'h3e;
		memory[16'h3bda] <= 8'h2a;
		memory[16'h3bdb] <= 8'h85;
		memory[16'h3bdc] <= 8'hbc;
		memory[16'h3bdd] <= 8'h9a;
		memory[16'h3bde] <= 8'h96;
		memory[16'h3bdf] <= 8'ha4;
		memory[16'h3be0] <= 8'hc8;
		memory[16'h3be1] <= 8'h52;
		memory[16'h3be2] <= 8'h95;
		memory[16'h3be3] <= 8'hb1;
		memory[16'h3be4] <= 8'ha3;
		memory[16'h3be5] <= 8'h32;
		memory[16'h3be6] <= 8'h99;
		memory[16'h3be7] <= 8'h70;
		memory[16'h3be8] <= 8'hee;
		memory[16'h3be9] <= 8'h5a;
		memory[16'h3bea] <= 8'hd1;
		memory[16'h3beb] <= 8'h74;
		memory[16'h3bec] <= 8'h6e;
		memory[16'h3bed] <= 8'h1c;
		memory[16'h3bee] <= 8'h35;
		memory[16'h3bef] <= 8'h60;
		memory[16'h3bf0] <= 8'h88;
		memory[16'h3bf1] <= 8'h17;
		memory[16'h3bf2] <= 8'hfe;
		memory[16'h3bf3] <= 8'hab;
		memory[16'h3bf4] <= 8'h13;
		memory[16'h3bf5] <= 8'h8c;
		memory[16'h3bf6] <= 8'h68;
		memory[16'h3bf7] <= 8'hb0;
		memory[16'h3bf8] <= 8'hca;
		memory[16'h3bf9] <= 8'h92;
		memory[16'h3bfa] <= 8'h36;
		memory[16'h3bfb] <= 8'h87;
		memory[16'h3bfc] <= 8'h2c;
		memory[16'h3bfd] <= 8'hcc;
		memory[16'h3bfe] <= 8'h2b;
		memory[16'h3bff] <= 8'hf4;
		memory[16'h3c00] <= 8'h1e;
		memory[16'h3c01] <= 8'hc0;
		memory[16'h3c02] <= 8'ha5;
		memory[16'h3c03] <= 8'hc1;
		memory[16'h3c04] <= 8'hf2;
		memory[16'h3c05] <= 8'h3e;
		memory[16'h3c06] <= 8'h31;
		memory[16'h3c07] <= 8'he1;
		memory[16'h3c08] <= 8'h98;
		memory[16'h3c09] <= 8'h3;
		memory[16'h3c0a] <= 8'h55;
		memory[16'h3c0b] <= 8'h7;
		memory[16'h3c0c] <= 8'h1f;
		memory[16'h3c0d] <= 8'h8a;
		memory[16'h3c0e] <= 8'h67;
		memory[16'h3c0f] <= 8'ha7;
		memory[16'h3c10] <= 8'ha1;
		memory[16'h3c11] <= 8'h65;
		memory[16'h3c12] <= 8'h52;
		memory[16'h3c13] <= 8'hb5;
		memory[16'h3c14] <= 8'hf1;
		memory[16'h3c15] <= 8'hba;
		memory[16'h3c16] <= 8'h65;
		memory[16'h3c17] <= 8'hbc;
		memory[16'h3c18] <= 8'h4c;
		memory[16'h3c19] <= 8'h9b;
		memory[16'h3c1a] <= 8'h43;
		memory[16'h3c1b] <= 8'h78;
		memory[16'h3c1c] <= 8'h68;
		memory[16'h3c1d] <= 8'h6e;
		memory[16'h3c1e] <= 8'h6d;
		memory[16'h3c1f] <= 8'h86;
		memory[16'h3c20] <= 8'h2e;
		memory[16'h3c21] <= 8'h12;
		memory[16'h3c22] <= 8'h48;
		memory[16'h3c23] <= 8'h21;
		memory[16'h3c24] <= 8'h51;
		memory[16'h3c25] <= 8'h79;
		memory[16'h3c26] <= 8'h2;
		memory[16'h3c27] <= 8'he9;
		memory[16'h3c28] <= 8'h7c;
		memory[16'h3c29] <= 8'h57;
		memory[16'h3c2a] <= 8'hf0;
		memory[16'h3c2b] <= 8'h9c;
		memory[16'h3c2c] <= 8'he1;
		memory[16'h3c2d] <= 8'h58;
		memory[16'h3c2e] <= 8'h43;
		memory[16'h3c2f] <= 8'h83;
		memory[16'h3c30] <= 8'hbd;
		memory[16'h3c31] <= 8'h96;
		memory[16'h3c32] <= 8'h38;
		memory[16'h3c33] <= 8'haf;
		memory[16'h3c34] <= 8'h50;
		memory[16'h3c35] <= 8'h9d;
		memory[16'h3c36] <= 8'h6b;
		memory[16'h3c37] <= 8'h9d;
		memory[16'h3c38] <= 8'h39;
		memory[16'h3c39] <= 8'hae;
		memory[16'h3c3a] <= 8'h15;
		memory[16'h3c3b] <= 8'ha1;
		memory[16'h3c3c] <= 8'h1c;
		memory[16'h3c3d] <= 8'h82;
		memory[16'h3c3e] <= 8'h27;
		memory[16'h3c3f] <= 8'h4a;
		memory[16'h3c40] <= 8'h95;
		memory[16'h3c41] <= 8'h6f;
		memory[16'h3c42] <= 8'h6b;
		memory[16'h3c43] <= 8'he6;
		memory[16'h3c44] <= 8'he9;
		memory[16'h3c45] <= 8'h6d;
		memory[16'h3c46] <= 8'hcf;
		memory[16'h3c47] <= 8'h65;
		memory[16'h3c48] <= 8'hc4;
		memory[16'h3c49] <= 8'hc0;
		memory[16'h3c4a] <= 8'h1;
		memory[16'h3c4b] <= 8'ha6;
		memory[16'h3c4c] <= 8'h18;
		memory[16'h3c4d] <= 8'h45;
		memory[16'h3c4e] <= 8'h29;
		memory[16'h3c4f] <= 8'hd5;
		memory[16'h3c50] <= 8'hdb;
		memory[16'h3c51] <= 8'h61;
		memory[16'h3c52] <= 8'h84;
		memory[16'h3c53] <= 8'h2b;
		memory[16'h3c54] <= 8'hfe;
		memory[16'h3c55] <= 8'hef;
		memory[16'h3c56] <= 8'hc8;
		memory[16'h3c57] <= 8'h37;
		memory[16'h3c58] <= 8'h9d;
		memory[16'h3c59] <= 8'hde;
		memory[16'h3c5a] <= 8'hd8;
		memory[16'h3c5b] <= 8'hb9;
		memory[16'h3c5c] <= 8'h60;
		memory[16'h3c5d] <= 8'h0;
		memory[16'h3c5e] <= 8'h4;
		memory[16'h3c5f] <= 8'hf5;
		memory[16'h3c60] <= 8'h6f;
		memory[16'h3c61] <= 8'h6f;
		memory[16'h3c62] <= 8'hdb;
		memory[16'h3c63] <= 8'h58;
		memory[16'h3c64] <= 8'hdd;
		memory[16'h3c65] <= 8'hab;
		memory[16'h3c66] <= 8'hbe;
		memory[16'h3c67] <= 8'ha1;
		memory[16'h3c68] <= 8'h6b;
		memory[16'h3c69] <= 8'hbf;
		memory[16'h3c6a] <= 8'h47;
		memory[16'h3c6b] <= 8'h83;
		memory[16'h3c6c] <= 8'h4;
		memory[16'h3c6d] <= 8'h70;
		memory[16'h3c6e] <= 8'h58;
		memory[16'h3c6f] <= 8'hdf;
		memory[16'h3c70] <= 8'hd1;
		memory[16'h3c71] <= 8'hdd;
		memory[16'h3c72] <= 8'hb;
		memory[16'h3c73] <= 8'hd0;
		memory[16'h3c74] <= 8'hcc;
		memory[16'h3c75] <= 8'hd3;
		memory[16'h3c76] <= 8'h7;
		memory[16'h3c77] <= 8'h6a;
		memory[16'h3c78] <= 8'hb1;
		memory[16'h3c79] <= 8'he0;
		memory[16'h3c7a] <= 8'h23;
		memory[16'h3c7b] <= 8'h12;
		memory[16'h3c7c] <= 8'he0;
		memory[16'h3c7d] <= 8'h27;
		memory[16'h3c7e] <= 8'h7;
		memory[16'h3c7f] <= 8'h4f;
		memory[16'h3c80] <= 8'h97;
		memory[16'h3c81] <= 8'he3;
		memory[16'h3c82] <= 8'ha8;
		memory[16'h3c83] <= 8'h74;
		memory[16'h3c84] <= 8'h8e;
		memory[16'h3c85] <= 8'h66;
		memory[16'h3c86] <= 8'h15;
		memory[16'h3c87] <= 8'hf9;
		memory[16'h3c88] <= 8'h25;
		memory[16'h3c89] <= 8'h5d;
		memory[16'h3c8a] <= 8'h7c;
		memory[16'h3c8b] <= 8'h2a;
		memory[16'h3c8c] <= 8'hcd;
		memory[16'h3c8d] <= 8'hd4;
		memory[16'h3c8e] <= 8'h9;
		memory[16'h3c8f] <= 8'h9f;
		memory[16'h3c90] <= 8'hb1;
		memory[16'h3c91] <= 8'h14;
		memory[16'h3c92] <= 8'h6f;
		memory[16'h3c93] <= 8'h7e;
		memory[16'h3c94] <= 8'he8;
		memory[16'h3c95] <= 8'h76;
		memory[16'h3c96] <= 8'he8;
		memory[16'h3c97] <= 8'h99;
		memory[16'h3c98] <= 8'h56;
		memory[16'h3c99] <= 8'hb;
		memory[16'h3c9a] <= 8'hab;
		memory[16'h3c9b] <= 8'h36;
		memory[16'h3c9c] <= 8'h33;
		memory[16'h3c9d] <= 8'hb3;
		memory[16'h3c9e] <= 8'h86;
		memory[16'h3c9f] <= 8'hca;
		memory[16'h3ca0] <= 8'h96;
		memory[16'h3ca1] <= 8'h2e;
		memory[16'h3ca2] <= 8'h3e;
		memory[16'h3ca3] <= 8'h24;
		memory[16'h3ca4] <= 8'h94;
		memory[16'h3ca5] <= 8'h53;
		memory[16'h3ca6] <= 8'h1d;
		memory[16'h3ca7] <= 8'hb9;
		memory[16'h3ca8] <= 8'hb0;
		memory[16'h3ca9] <= 8'h99;
		memory[16'h3caa] <= 8'he3;
		memory[16'h3cab] <= 8'h7e;
		memory[16'h3cac] <= 8'h6d;
		memory[16'h3cad] <= 8'hed;
		memory[16'h3cae] <= 8'h1d;
		memory[16'h3caf] <= 8'h1f;
		memory[16'h3cb0] <= 8'h1;
		memory[16'h3cb1] <= 8'h8c;
		memory[16'h3cb2] <= 8'h9d;
		memory[16'h3cb3] <= 8'he9;
		memory[16'h3cb4] <= 8'h2;
		memory[16'h3cb5] <= 8'h85;
		memory[16'h3cb6] <= 8'h83;
		memory[16'h3cb7] <= 8'h59;
		memory[16'h3cb8] <= 8'h90;
		memory[16'h3cb9] <= 8'h2e;
		memory[16'h3cba] <= 8'h8f;
		memory[16'h3cbb] <= 8'hc3;
		memory[16'h3cbc] <= 8'he1;
		memory[16'h3cbd] <= 8'h15;
		memory[16'h3cbe] <= 8'h8d;
		memory[16'h3cbf] <= 8'h77;
		memory[16'h3cc0] <= 8'h43;
		memory[16'h3cc1] <= 8'hcb;
		memory[16'h3cc2] <= 8'h9b;
		memory[16'h3cc3] <= 8'hd7;
		memory[16'h3cc4] <= 8'h1f;
		memory[16'h3cc5] <= 8'hb8;
		memory[16'h3cc6] <= 8'h91;
		memory[16'h3cc7] <= 8'hcf;
		memory[16'h3cc8] <= 8'h51;
		memory[16'h3cc9] <= 8'h74;
		memory[16'h3cca] <= 8'h4d;
		memory[16'h3ccb] <= 8'hbf;
		memory[16'h3ccc] <= 8'h61;
		memory[16'h3ccd] <= 8'h6a;
		memory[16'h3cce] <= 8'hde;
		memory[16'h3ccf] <= 8'h63;
		memory[16'h3cd0] <= 8'hf6;
		memory[16'h3cd1] <= 8'h7b;
		memory[16'h3cd2] <= 8'h4c;
		memory[16'h3cd3] <= 8'hf9;
		memory[16'h3cd4] <= 8'h0;
		memory[16'h3cd5] <= 8'hcf;
		memory[16'h3cd6] <= 8'h52;
		memory[16'h3cd7] <= 8'h90;
		memory[16'h3cd8] <= 8'hfe;
		memory[16'h3cd9] <= 8'he1;
		memory[16'h3cda] <= 8'h54;
		memory[16'h3cdb] <= 8'hdf;
		memory[16'h3cdc] <= 8'hf7;
		memory[16'h3cdd] <= 8'he1;
		memory[16'h3cde] <= 8'h57;
		memory[16'h3cdf] <= 8'h3a;
		memory[16'h3ce0] <= 8'had;
		memory[16'h3ce1] <= 8'hf2;
		memory[16'h3ce2] <= 8'h12;
		memory[16'h3ce3] <= 8'hcc;
		memory[16'h3ce4] <= 8'hab;
		memory[16'h3ce5] <= 8'ha3;
		memory[16'h3ce6] <= 8'h9b;
		memory[16'h3ce7] <= 8'hfc;
		memory[16'h3ce8] <= 8'h17;
		memory[16'h3ce9] <= 8'he9;
		memory[16'h3cea] <= 8'hbb;
		memory[16'h3ceb] <= 8'h79;
		memory[16'h3cec] <= 8'h53;
		memory[16'h3ced] <= 8'h99;
		memory[16'h3cee] <= 8'hdc;
		memory[16'h3cef] <= 8'h4a;
		memory[16'h3cf0] <= 8'h14;
		memory[16'h3cf1] <= 8'h28;
		memory[16'h3cf2] <= 8'h43;
		memory[16'h3cf3] <= 8'h14;
		memory[16'h3cf4] <= 8'hf8;
		memory[16'h3cf5] <= 8'h95;
		memory[16'h3cf6] <= 8'ha5;
		memory[16'h3cf7] <= 8'hf6;
		memory[16'h3cf8] <= 8'h76;
		memory[16'h3cf9] <= 8'hf9;
		memory[16'h3cfa] <= 8'hd5;
		memory[16'h3cfb] <= 8'h6d;
		memory[16'h3cfc] <= 8'hda;
		memory[16'h3cfd] <= 8'h2c;
		memory[16'h3cfe] <= 8'ha8;
		memory[16'h3cff] <= 8'h87;
		memory[16'h3d00] <= 8'h1f;
		memory[16'h3d01] <= 8'hba;
		memory[16'h3d02] <= 8'h53;
		memory[16'h3d03] <= 8'hca;
		memory[16'h3d04] <= 8'h5d;
		memory[16'h3d05] <= 8'hef;
		memory[16'h3d06] <= 8'hc6;
		memory[16'h3d07] <= 8'h74;
		memory[16'h3d08] <= 8'hd8;
		memory[16'h3d09] <= 8'h82;
		memory[16'h3d0a] <= 8'hed;
		memory[16'h3d0b] <= 8'h2b;
		memory[16'h3d0c] <= 8'h1b;
		memory[16'h3d0d] <= 8'hc9;
		memory[16'h3d0e] <= 8'h75;
		memory[16'h3d0f] <= 8'h30;
		memory[16'h3d10] <= 8'hf2;
		memory[16'h3d11] <= 8'hb8;
		memory[16'h3d12] <= 8'h44;
		memory[16'h3d13] <= 8'hea;
		memory[16'h3d14] <= 8'h4d;
		memory[16'h3d15] <= 8'he9;
		memory[16'h3d16] <= 8'he0;
		memory[16'h3d17] <= 8'hc4;
		memory[16'h3d18] <= 8'he2;
		memory[16'h3d19] <= 8'hb5;
		memory[16'h3d1a] <= 8'h31;
		memory[16'h3d1b] <= 8'hbd;
		memory[16'h3d1c] <= 8'he2;
		memory[16'h3d1d] <= 8'hd9;
		memory[16'h3d1e] <= 8'h44;
		memory[16'h3d1f] <= 8'h1;
		memory[16'h3d20] <= 8'h93;
		memory[16'h3d21] <= 8'h98;
		memory[16'h3d22] <= 8'hcb;
		memory[16'h3d23] <= 8'hf0;
		memory[16'h3d24] <= 8'h87;
		memory[16'h3d25] <= 8'h91;
		memory[16'h3d26] <= 8'h65;
		memory[16'h3d27] <= 8'h5f;
		memory[16'h3d28] <= 8'h13;
		memory[16'h3d29] <= 8'h52;
		memory[16'h3d2a] <= 8'h8a;
		memory[16'h3d2b] <= 8'h2f;
		memory[16'h3d2c] <= 8'h1c;
		memory[16'h3d2d] <= 8'h0;
		memory[16'h3d2e] <= 8'h5f;
		memory[16'h3d2f] <= 8'he;
		memory[16'h3d30] <= 8'hb8;
		memory[16'h3d31] <= 8'ha3;
		memory[16'h3d32] <= 8'hf8;
		memory[16'h3d33] <= 8'h6;
		memory[16'h3d34] <= 8'h8d;
		memory[16'h3d35] <= 8'hd8;
		memory[16'h3d36] <= 8'hca;
		memory[16'h3d37] <= 8'h6f;
		memory[16'h3d38] <= 8'h8d;
		memory[16'h3d39] <= 8'hfb;
		memory[16'h3d3a] <= 8'h2c;
		memory[16'h3d3b] <= 8'h6f;
		memory[16'h3d3c] <= 8'hd5;
		memory[16'h3d3d] <= 8'h71;
		memory[16'h3d3e] <= 8'h70;
		memory[16'h3d3f] <= 8'h68;
		memory[16'h3d40] <= 8'h9;
		memory[16'h3d41] <= 8'h3b;
		memory[16'h3d42] <= 8'h59;
		memory[16'h3d43] <= 8'h90;
		memory[16'h3d44] <= 8'hcd;
		memory[16'h3d45] <= 8'hbe;
		memory[16'h3d46] <= 8'hef;
		memory[16'h3d47] <= 8'he0;
		memory[16'h3d48] <= 8'h10;
		memory[16'h3d49] <= 8'h79;
		memory[16'h3d4a] <= 8'hf;
		memory[16'h3d4b] <= 8'h2c;
		memory[16'h3d4c] <= 8'h79;
		memory[16'h3d4d] <= 8'h6e;
		memory[16'h3d4e] <= 8'h3a;
		memory[16'h3d4f] <= 8'h32;
		memory[16'h3d50] <= 8'h12;
		memory[16'h3d51] <= 8'h32;
		memory[16'h3d52] <= 8'h38;
		memory[16'h3d53] <= 8'h9f;
		memory[16'h3d54] <= 8'ha;
		memory[16'h3d55] <= 8'h2;
		memory[16'h3d56] <= 8'he;
		memory[16'h3d57] <= 8'h98;
		memory[16'h3d58] <= 8'hfd;
		memory[16'h3d59] <= 8'h3b;
		memory[16'h3d5a] <= 8'h7;
		memory[16'h3d5b] <= 8'hd2;
		memory[16'h3d5c] <= 8'hac;
		memory[16'h3d5d] <= 8'h78;
		memory[16'h3d5e] <= 8'h3b;
		memory[16'h3d5f] <= 8'hb5;
		memory[16'h3d60] <= 8'hb3;
		memory[16'h3d61] <= 8'h94;
		memory[16'h3d62] <= 8'h45;
		memory[16'h3d63] <= 8'h80;
		memory[16'h3d64] <= 8'h52;
		memory[16'h3d65] <= 8'h34;
		memory[16'h3d66] <= 8'h61;
		memory[16'h3d67] <= 8'h62;
		memory[16'h3d68] <= 8'had;
		memory[16'h3d69] <= 8'h70;
		memory[16'h3d6a] <= 8'h8f;
		memory[16'h3d6b] <= 8'h27;
		memory[16'h3d6c] <= 8'hdf;
		memory[16'h3d6d] <= 8'hc9;
		memory[16'h3d6e] <= 8'h59;
		memory[16'h3d6f] <= 8'hf1;
		memory[16'h3d70] <= 8'hfc;
		memory[16'h3d71] <= 8'h91;
		memory[16'h3d72] <= 8'h90;
		memory[16'h3d73] <= 8'h6;
		memory[16'h3d74] <= 8'h93;
		memory[16'h3d75] <= 8'h9e;
		memory[16'h3d76] <= 8'h9e;
		memory[16'h3d77] <= 8'h90;
		memory[16'h3d78] <= 8'hd9;
		memory[16'h3d79] <= 8'ha6;
		memory[16'h3d7a] <= 8'h63;
		memory[16'h3d7b] <= 8'h85;
		memory[16'h3d7c] <= 8'h1e;
		memory[16'h3d7d] <= 8'h9e;
		memory[16'h3d7e] <= 8'h3a;
		memory[16'h3d7f] <= 8'hd1;
		memory[16'h3d80] <= 8'h32;
		memory[16'h3d81] <= 8'h7f;
		memory[16'h3d82] <= 8'h52;
		memory[16'h3d83] <= 8'h84;
		memory[16'h3d84] <= 8'hb3;
		memory[16'h3d85] <= 8'hb3;
		memory[16'h3d86] <= 8'he6;
		memory[16'h3d87] <= 8'h61;
		memory[16'h3d88] <= 8'h23;
		memory[16'h3d89] <= 8'h75;
		memory[16'h3d8a] <= 8'h88;
		memory[16'h3d8b] <= 8'h2;
		memory[16'h3d8c] <= 8'h3f;
		memory[16'h3d8d] <= 8'he1;
		memory[16'h3d8e] <= 8'hf3;
		memory[16'h3d8f] <= 8'h3b;
		memory[16'h3d90] <= 8'h72;
		memory[16'h3d91] <= 8'h83;
		memory[16'h3d92] <= 8'h41;
		memory[16'h3d93] <= 8'h5;
		memory[16'h3d94] <= 8'h22;
		memory[16'h3d95] <= 8'he0;
		memory[16'h3d96] <= 8'h95;
		memory[16'h3d97] <= 8'hfb;
		memory[16'h3d98] <= 8'h86;
		memory[16'h3d99] <= 8'hf8;
		memory[16'h3d9a] <= 8'h81;
		memory[16'h3d9b] <= 8'ha4;
		memory[16'h3d9c] <= 8'h96;
		memory[16'h3d9d] <= 8'hbb;
		memory[16'h3d9e] <= 8'h75;
		memory[16'h3d9f] <= 8'hc8;
		memory[16'h3da0] <= 8'h3b;
		memory[16'h3da1] <= 8'hc7;
		memory[16'h3da2] <= 8'h4c;
		memory[16'h3da3] <= 8'hee;
		memory[16'h3da4] <= 8'h7a;
		memory[16'h3da5] <= 8'h33;
		memory[16'h3da6] <= 8'h4f;
		memory[16'h3da7] <= 8'h9e;
		memory[16'h3da8] <= 8'ha8;
		memory[16'h3da9] <= 8'hd7;
		memory[16'h3daa] <= 8'ha0;
		memory[16'h3dab] <= 8'he7;
		memory[16'h3dac] <= 8'hb8;
		memory[16'h3dad] <= 8'h94;
		memory[16'h3dae] <= 8'h22;
		memory[16'h3daf] <= 8'h2a;
		memory[16'h3db0] <= 8'h17;
		memory[16'h3db1] <= 8'h64;
		memory[16'h3db2] <= 8'h2f;
		memory[16'h3db3] <= 8'h39;
		memory[16'h3db4] <= 8'h44;
		memory[16'h3db5] <= 8'hc5;
		memory[16'h3db6] <= 8'h35;
		memory[16'h3db7] <= 8'hca;
		memory[16'h3db8] <= 8'hbd;
		memory[16'h3db9] <= 8'hb6;
		memory[16'h3dba] <= 8'h6e;
		memory[16'h3dbb] <= 8'h54;
		memory[16'h3dbc] <= 8'h71;
		memory[16'h3dbd] <= 8'he3;
		memory[16'h3dbe] <= 8'h1c;
		memory[16'h3dbf] <= 8'hac;
		memory[16'h3dc0] <= 8'hab;
		memory[16'h3dc1] <= 8'h69;
		memory[16'h3dc2] <= 8'h9b;
		memory[16'h3dc3] <= 8'h25;
		memory[16'h3dc4] <= 8'h9c;
		memory[16'h3dc5] <= 8'hea;
		memory[16'h3dc6] <= 8'hc3;
		memory[16'h3dc7] <= 8'h44;
		memory[16'h3dc8] <= 8'hc2;
		memory[16'h3dc9] <= 8'h64;
		memory[16'h3dca] <= 8'h2c;
		memory[16'h3dcb] <= 8'h7a;
		memory[16'h3dcc] <= 8'hf8;
		memory[16'h3dcd] <= 8'h4e;
		memory[16'h3dce] <= 8'ha5;
		memory[16'h3dcf] <= 8'hf;
		memory[16'h3dd0] <= 8'hb2;
		memory[16'h3dd1] <= 8'hd4;
		memory[16'h3dd2] <= 8'h49;
		memory[16'h3dd3] <= 8'hf6;
		memory[16'h3dd4] <= 8'h99;
		memory[16'h3dd5] <= 8'h7e;
		memory[16'h3dd6] <= 8'hc0;
		memory[16'h3dd7] <= 8'h57;
		memory[16'h3dd8] <= 8'h34;
		memory[16'h3dd9] <= 8'h2e;
		memory[16'h3dda] <= 8'hab;
		memory[16'h3ddb] <= 8'ha5;
		memory[16'h3ddc] <= 8'h12;
		memory[16'h3ddd] <= 8'hc7;
		memory[16'h3dde] <= 8'h52;
		memory[16'h3ddf] <= 8'hbd;
		memory[16'h3de0] <= 8'h30;
		memory[16'h3de1] <= 8'hed;
		memory[16'h3de2] <= 8'he2;
		memory[16'h3de3] <= 8'hcc;
		memory[16'h3de4] <= 8'hd7;
		memory[16'h3de5] <= 8'ha6;
		memory[16'h3de6] <= 8'h11;
		memory[16'h3de7] <= 8'h99;
		memory[16'h3de8] <= 8'ha;
		memory[16'h3de9] <= 8'h3d;
		memory[16'h3dea] <= 8'h14;
		memory[16'h3deb] <= 8'h2;
		memory[16'h3dec] <= 8'h8b;
		memory[16'h3ded] <= 8'hb9;
		memory[16'h3dee] <= 8'h11;
		memory[16'h3def] <= 8'h3e;
		memory[16'h3df0] <= 8'h8d;
		memory[16'h3df1] <= 8'h5a;
		memory[16'h3df2] <= 8'h34;
		memory[16'h3df3] <= 8'h27;
		memory[16'h3df4] <= 8'hd8;
		memory[16'h3df5] <= 8'hf5;
		memory[16'h3df6] <= 8'h7e;
		memory[16'h3df7] <= 8'hc;
		memory[16'h3df8] <= 8'h23;
		memory[16'h3df9] <= 8'h29;
		memory[16'h3dfa] <= 8'hb2;
		memory[16'h3dfb] <= 8'h35;
		memory[16'h3dfc] <= 8'hf0;
		memory[16'h3dfd] <= 8'h4;
		memory[16'h3dfe] <= 8'hf2;
		memory[16'h3dff] <= 8'h21;
		memory[16'h3e00] <= 8'hf1;
		memory[16'h3e01] <= 8'hd5;
		memory[16'h3e02] <= 8'hed;
		memory[16'h3e03] <= 8'hc8;
		memory[16'h3e04] <= 8'h7b;
		memory[16'h3e05] <= 8'hfe;
		memory[16'h3e06] <= 8'h62;
		memory[16'h3e07] <= 8'h85;
		memory[16'h3e08] <= 8'h3b;
		memory[16'h3e09] <= 8'h76;
		memory[16'h3e0a] <= 8'h87;
		memory[16'h3e0b] <= 8'hc7;
		memory[16'h3e0c] <= 8'h2f;
		memory[16'h3e0d] <= 8'h98;
		memory[16'h3e0e] <= 8'h5;
		memory[16'h3e0f] <= 8'hbc;
		memory[16'h3e10] <= 8'hf3;
		memory[16'h3e11] <= 8'h39;
		memory[16'h3e12] <= 8'he3;
		memory[16'h3e13] <= 8'hcb;
		memory[16'h3e14] <= 8'h2e;
		memory[16'h3e15] <= 8'h61;
		memory[16'h3e16] <= 8'hd8;
		memory[16'h3e17] <= 8'h52;
		memory[16'h3e18] <= 8'h8a;
		memory[16'h3e19] <= 8'h8a;
		memory[16'h3e1a] <= 8'h87;
		memory[16'h3e1b] <= 8'h7b;
		memory[16'h3e1c] <= 8'h8e;
		memory[16'h3e1d] <= 8'h7a;
		memory[16'h3e1e] <= 8'h9c;
		memory[16'h3e1f] <= 8'h7f;
		memory[16'h3e20] <= 8'h4f;
		memory[16'h3e21] <= 8'h89;
		memory[16'h3e22] <= 8'h47;
		memory[16'h3e23] <= 8'hca;
		memory[16'h3e24] <= 8'h88;
		memory[16'h3e25] <= 8'ha9;
		memory[16'h3e26] <= 8'h4f;
		memory[16'h3e27] <= 8'hc3;
		memory[16'h3e28] <= 8'h1f;
		memory[16'h3e29] <= 8'hd6;
		memory[16'h3e2a] <= 8'h8a;
		memory[16'h3e2b] <= 8'h4e;
		memory[16'h3e2c] <= 8'h6e;
		memory[16'h3e2d] <= 8'h8f;
		memory[16'h3e2e] <= 8'hb;
		memory[16'h3e2f] <= 8'h61;
		memory[16'h3e30] <= 8'hc9;
		memory[16'h3e31] <= 8'hee;
		memory[16'h3e32] <= 8'h2d;
		memory[16'h3e33] <= 8'hf7;
		memory[16'h3e34] <= 8'h50;
		memory[16'h3e35] <= 8'h5;
		memory[16'h3e36] <= 8'h49;
		memory[16'h3e37] <= 8'hda;
		memory[16'h3e38] <= 8'h8f;
		memory[16'h3e39] <= 8'hd1;
		memory[16'h3e3a] <= 8'h55;
		memory[16'h3e3b] <= 8'h1d;
		memory[16'h3e3c] <= 8'h4b;
		memory[16'h3e3d] <= 8'hf1;
		memory[16'h3e3e] <= 8'h9c;
		memory[16'h3e3f] <= 8'h9a;
		memory[16'h3e40] <= 8'h7b;
		memory[16'h3e41] <= 8'he3;
		memory[16'h3e42] <= 8'h64;
		memory[16'h3e43] <= 8'h3;
		memory[16'h3e44] <= 8'h8d;
		memory[16'h3e45] <= 8'hb3;
		memory[16'h3e46] <= 8'hc6;
		memory[16'h3e47] <= 8'hac;
		memory[16'h3e48] <= 8'h89;
		memory[16'h3e49] <= 8'h51;
		memory[16'h3e4a] <= 8'hfb;
		memory[16'h3e4b] <= 8'hf7;
		memory[16'h3e4c] <= 8'he0;
		memory[16'h3e4d] <= 8'h6;
		memory[16'h3e4e] <= 8'h59;
		memory[16'h3e4f] <= 8'ha9;
		memory[16'h3e50] <= 8'hf4;
		memory[16'h3e51] <= 8'h86;
		memory[16'h3e52] <= 8'ha1;
		memory[16'h3e53] <= 8'h44;
		memory[16'h3e54] <= 8'h8b;
		memory[16'h3e55] <= 8'hea;
		memory[16'h3e56] <= 8'h1f;
		memory[16'h3e57] <= 8'h1a;
		memory[16'h3e58] <= 8'hbb;
		memory[16'h3e59] <= 8'h74;
		memory[16'h3e5a] <= 8'h37;
		memory[16'h3e5b] <= 8'h6;
		memory[16'h3e5c] <= 8'h66;
		memory[16'h3e5d] <= 8'hd3;
		memory[16'h3e5e] <= 8'ha0;
		memory[16'h3e5f] <= 8'he1;
		memory[16'h3e60] <= 8'hb6;
		memory[16'h3e61] <= 8'h4;
		memory[16'h3e62] <= 8'he4;
		memory[16'h3e63] <= 8'h43;
		memory[16'h3e64] <= 8'hb7;
		memory[16'h3e65] <= 8'haa;
		memory[16'h3e66] <= 8'hf0;
		memory[16'h3e67] <= 8'h40;
		memory[16'h3e68] <= 8'hfb;
		memory[16'h3e69] <= 8'heb;
		memory[16'h3e6a] <= 8'h38;
		memory[16'h3e6b] <= 8'hdc;
		memory[16'h3e6c] <= 8'hf1;
		memory[16'h3e6d] <= 8'h91;
		memory[16'h3e6e] <= 8'h85;
		memory[16'h3e6f] <= 8'he5;
		memory[16'h3e70] <= 8'h17;
		memory[16'h3e71] <= 8'h26;
		memory[16'h3e72] <= 8'h2a;
		memory[16'h3e73] <= 8'ha2;
		memory[16'h3e74] <= 8'h11;
		memory[16'h3e75] <= 8'h49;
		memory[16'h3e76] <= 8'hbc;
		memory[16'h3e77] <= 8'hcc;
		memory[16'h3e78] <= 8'hbd;
		memory[16'h3e79] <= 8'hf3;
		memory[16'h3e7a] <= 8'hd3;
		memory[16'h3e7b] <= 8'h23;
		memory[16'h3e7c] <= 8'hc6;
		memory[16'h3e7d] <= 8'h73;
		memory[16'h3e7e] <= 8'h4;
		memory[16'h3e7f] <= 8'h7c;
		memory[16'h3e80] <= 8'h78;
		memory[16'h3e81] <= 8'he8;
		memory[16'h3e82] <= 8'hc0;
		memory[16'h3e83] <= 8'h2f;
		memory[16'h3e84] <= 8'h93;
		memory[16'h3e85] <= 8'hb0;
		memory[16'h3e86] <= 8'h70;
		memory[16'h3e87] <= 8'h8e;
		memory[16'h3e88] <= 8'h9b;
		memory[16'h3e89] <= 8'ha8;
		memory[16'h3e8a] <= 8'h6a;
		memory[16'h3e8b] <= 8'h8c;
		memory[16'h3e8c] <= 8'h39;
		memory[16'h3e8d] <= 8'hf0;
		memory[16'h3e8e] <= 8'h71;
		memory[16'h3e8f] <= 8'h50;
		memory[16'h3e90] <= 8'h16;
		memory[16'h3e91] <= 8'h9b;
		memory[16'h3e92] <= 8'hf2;
		memory[16'h3e93] <= 8'h27;
		memory[16'h3e94] <= 8'he4;
		memory[16'h3e95] <= 8'hae;
		memory[16'h3e96] <= 8'hf4;
		memory[16'h3e97] <= 8'ha2;
		memory[16'h3e98] <= 8'ha1;
		memory[16'h3e99] <= 8'hc7;
		memory[16'h3e9a] <= 8'hc5;
		memory[16'h3e9b] <= 8'h67;
		memory[16'h3e9c] <= 8'h3a;
		memory[16'h3e9d] <= 8'hca;
		memory[16'h3e9e] <= 8'he3;
		memory[16'h3e9f] <= 8'hb2;
		memory[16'h3ea0] <= 8'hb2;
		memory[16'h3ea1] <= 8'ha3;
		memory[16'h3ea2] <= 8'he2;
		memory[16'h3ea3] <= 8'h45;
		memory[16'h3ea4] <= 8'h53;
		memory[16'h3ea5] <= 8'h52;
		memory[16'h3ea6] <= 8'hd4;
		memory[16'h3ea7] <= 8'hee;
		memory[16'h3ea8] <= 8'hfa;
		memory[16'h3ea9] <= 8'h3e;
		memory[16'h3eaa] <= 8'h7a;
		memory[16'h3eab] <= 8'h33;
		memory[16'h3eac] <= 8'h2e;
		memory[16'h3ead] <= 8'hec;
		memory[16'h3eae] <= 8'h83;
		memory[16'h3eaf] <= 8'h45;
		memory[16'h3eb0] <= 8'h87;
		memory[16'h3eb1] <= 8'h75;
		memory[16'h3eb2] <= 8'h6c;
		memory[16'h3eb3] <= 8'h6c;
		memory[16'h3eb4] <= 8'h23;
		memory[16'h3eb5] <= 8'h60;
		memory[16'h3eb6] <= 8'he;
		memory[16'h3eb7] <= 8'hc4;
		memory[16'h3eb8] <= 8'h27;
		memory[16'h3eb9] <= 8'hd3;
		memory[16'h3eba] <= 8'h2b;
		memory[16'h3ebb] <= 8'h62;
		memory[16'h3ebc] <= 8'h9d;
		memory[16'h3ebd] <= 8'he;
		memory[16'h3ebe] <= 8'h14;
		memory[16'h3ebf] <= 8'h50;
		memory[16'h3ec0] <= 8'hb2;
		memory[16'h3ec1] <= 8'hf6;
		memory[16'h3ec2] <= 8'h95;
		memory[16'h3ec3] <= 8'h5;
		memory[16'h3ec4] <= 8'h48;
		memory[16'h3ec5] <= 8'h69;
		memory[16'h3ec6] <= 8'hf4;
		memory[16'h3ec7] <= 8'h42;
		memory[16'h3ec8] <= 8'ha8;
		memory[16'h3ec9] <= 8'h6e;
		memory[16'h3eca] <= 8'h75;
		memory[16'h3ecb] <= 8'hd6;
		memory[16'h3ecc] <= 8'h5a;
		memory[16'h3ecd] <= 8'hf8;
		memory[16'h3ece] <= 8'h1b;
		memory[16'h3ecf] <= 8'he2;
		memory[16'h3ed0] <= 8'h6d;
		memory[16'h3ed1] <= 8'h88;
		memory[16'h3ed2] <= 8'h4e;
		memory[16'h3ed3] <= 8'h90;
		memory[16'h3ed4] <= 8'he8;
		memory[16'h3ed5] <= 8'h5c;
		memory[16'h3ed6] <= 8'h54;
		memory[16'h3ed7] <= 8'h10;
		memory[16'h3ed8] <= 8'h2f;
		memory[16'h3ed9] <= 8'h7f;
		memory[16'h3eda] <= 8'h72;
		memory[16'h3edb] <= 8'hcd;
		memory[16'h3edc] <= 8'h8e;
		memory[16'h3edd] <= 8'h86;
		memory[16'h3ede] <= 8'h1d;
		memory[16'h3edf] <= 8'h40;
		memory[16'h3ee0] <= 8'h7d;
		memory[16'h3ee1] <= 8'hb2;
		memory[16'h3ee2] <= 8'h45;
		memory[16'h3ee3] <= 8'hc5;
		memory[16'h3ee4] <= 8'h1c;
		memory[16'h3ee5] <= 8'h39;
		memory[16'h3ee6] <= 8'h8;
		memory[16'h3ee7] <= 8'hc4;
		memory[16'h3ee8] <= 8'ha8;
		memory[16'h3ee9] <= 8'h7d;
		memory[16'h3eea] <= 8'h9a;
		memory[16'h3eeb] <= 8'h2;
		memory[16'h3eec] <= 8'h76;
		memory[16'h3eed] <= 8'hb6;
		memory[16'h3eee] <= 8'he4;
		memory[16'h3eef] <= 8'he3;
		memory[16'h3ef0] <= 8'h3e;
		memory[16'h3ef1] <= 8'h32;
		memory[16'h3ef2] <= 8'h74;
		memory[16'h3ef3] <= 8'h26;
		memory[16'h3ef4] <= 8'h8e;
		memory[16'h3ef5] <= 8'hc8;
		memory[16'h3ef6] <= 8'h36;
		memory[16'h3ef7] <= 8'hbe;
		memory[16'h3ef8] <= 8'h48;
		memory[16'h3ef9] <= 8'ha8;
		memory[16'h3efa] <= 8'h8b;
		memory[16'h3efb] <= 8'hd6;
		memory[16'h3efc] <= 8'h2f;
		memory[16'h3efd] <= 8'ha8;
		memory[16'h3efe] <= 8'h16;
		memory[16'h3eff] <= 8'hac;
		memory[16'h3f00] <= 8'h5a;
		memory[16'h3f01] <= 8'h5b;
		memory[16'h3f02] <= 8'h71;
		memory[16'h3f03] <= 8'h76;
		memory[16'h3f04] <= 8'h95;
		memory[16'h3f05] <= 8'h79;
		memory[16'h3f06] <= 8'h3a;
		memory[16'h3f07] <= 8'h3d;
		memory[16'h3f08] <= 8'hf7;
		memory[16'h3f09] <= 8'hd5;
		memory[16'h3f0a] <= 8'h3f;
		memory[16'h3f0b] <= 8'h6d;
		memory[16'h3f0c] <= 8'h8b;
		memory[16'h3f0d] <= 8'h24;
		memory[16'h3f0e] <= 8'h50;
		memory[16'h3f0f] <= 8'hc9;
		memory[16'h3f10] <= 8'h56;
		memory[16'h3f11] <= 8'hc4;
		memory[16'h3f12] <= 8'hef;
		memory[16'h3f13] <= 8'he5;
		memory[16'h3f14] <= 8'h8d;
		memory[16'h3f15] <= 8'h26;
		memory[16'h3f16] <= 8'ha3;
		memory[16'h3f17] <= 8'hd5;
		memory[16'h3f18] <= 8'hce;
		memory[16'h3f19] <= 8'h2e;
		memory[16'h3f1a] <= 8'hab;
		memory[16'h3f1b] <= 8'hfd;
		memory[16'h3f1c] <= 8'hd6;
		memory[16'h3f1d] <= 8'hc1;
		memory[16'h3f1e] <= 8'ha9;
		memory[16'h3f1f] <= 8'h30;
		memory[16'h3f20] <= 8'h1c;
		memory[16'h3f21] <= 8'h1b;
		memory[16'h3f22] <= 8'ha7;
		memory[16'h3f23] <= 8'hb1;
		memory[16'h3f24] <= 8'h94;
		memory[16'h3f25] <= 8'he1;
		memory[16'h3f26] <= 8'hee;
		memory[16'h3f27] <= 8'h8b;
		memory[16'h3f28] <= 8'hb6;
		memory[16'h3f29] <= 8'h2e;
		memory[16'h3f2a] <= 8'hf8;
		memory[16'h3f2b] <= 8'h41;
		memory[16'h3f2c] <= 8'h52;
		memory[16'h3f2d] <= 8'h49;
		memory[16'h3f2e] <= 8'ha;
		memory[16'h3f2f] <= 8'ha8;
		memory[16'h3f30] <= 8'hd;
		memory[16'h3f31] <= 8'hfa;
		memory[16'h3f32] <= 8'h8d;
		memory[16'h3f33] <= 8'h9a;
		memory[16'h3f34] <= 8'h20;
		memory[16'h3f35] <= 8'h30;
		memory[16'h3f36] <= 8'h6f;
		memory[16'h3f37] <= 8'hee;
		memory[16'h3f38] <= 8'h5e;
		memory[16'h3f39] <= 8'h1a;
		memory[16'h3f3a] <= 8'hec;
		memory[16'h3f3b] <= 8'h34;
		memory[16'h3f3c] <= 8'hdb;
		memory[16'h3f3d] <= 8'h95;
		memory[16'h3f3e] <= 8'h65;
		memory[16'h3f3f] <= 8'hf8;
		memory[16'h3f40] <= 8'hb0;
		memory[16'h3f41] <= 8'hc;
		memory[16'h3f42] <= 8'ha9;
		memory[16'h3f43] <= 8'h45;
		memory[16'h3f44] <= 8'hed;
		memory[16'h3f45] <= 8'h98;
		memory[16'h3f46] <= 8'hd0;
		memory[16'h3f47] <= 8'ha4;
		memory[16'h3f48] <= 8'hc6;
		memory[16'h3f49] <= 8'hc9;
		memory[16'h3f4a] <= 8'he5;
		memory[16'h3f4b] <= 8'h18;
		memory[16'h3f4c] <= 8'h12;
		memory[16'h3f4d] <= 8'hf0;
		memory[16'h3f4e] <= 8'hc0;
		memory[16'h3f4f] <= 8'h1f;
		memory[16'h3f50] <= 8'hea;
		memory[16'h3f51] <= 8'h4e;
		memory[16'h3f52] <= 8'hba;
		memory[16'h3f53] <= 8'ha;
		memory[16'h3f54] <= 8'h7e;
		memory[16'h3f55] <= 8'h29;
		memory[16'h3f56] <= 8'hf8;
		memory[16'h3f57] <= 8'hdd;
		memory[16'h3f58] <= 8'h44;
		memory[16'h3f59] <= 8'he4;
		memory[16'h3f5a] <= 8'h11;
		memory[16'h3f5b] <= 8'h1f;
		memory[16'h3f5c] <= 8'h7a;
		memory[16'h3f5d] <= 8'h76;
		memory[16'h3f5e] <= 8'h17;
		memory[16'h3f5f] <= 8'h2a;
		memory[16'h3f60] <= 8'h82;
		memory[16'h3f61] <= 8'hc1;
		memory[16'h3f62] <= 8'h6f;
		memory[16'h3f63] <= 8'h70;
		memory[16'h3f64] <= 8'h59;
		memory[16'h3f65] <= 8'h40;
		memory[16'h3f66] <= 8'h14;
		memory[16'h3f67] <= 8'h1f;
		memory[16'h3f68] <= 8'h9;
		memory[16'h3f69] <= 8'hf9;
		memory[16'h3f6a] <= 8'h37;
		memory[16'h3f6b] <= 8'h1b;
		memory[16'h3f6c] <= 8'he9;
		memory[16'h3f6d] <= 8'hf7;
		memory[16'h3f6e] <= 8'h3a;
		memory[16'h3f6f] <= 8'hd3;
		memory[16'h3f70] <= 8'h45;
		memory[16'h3f71] <= 8'hf4;
		memory[16'h3f72] <= 8'hdd;
		memory[16'h3f73] <= 8'hc4;
		memory[16'h3f74] <= 8'h1e;
		memory[16'h3f75] <= 8'hd6;
		memory[16'h3f76] <= 8'ha1;
		memory[16'h3f77] <= 8'h62;
		memory[16'h3f78] <= 8'hba;
		memory[16'h3f79] <= 8'hb2;
		memory[16'h3f7a] <= 8'h81;
		memory[16'h3f7b] <= 8'h34;
		memory[16'h3f7c] <= 8'h29;
		memory[16'h3f7d] <= 8'h99;
		memory[16'h3f7e] <= 8'h5f;
		memory[16'h3f7f] <= 8'hab;
		memory[16'h3f80] <= 8'h5a;
		memory[16'h3f81] <= 8'hce;
		memory[16'h3f82] <= 8'h1b;
		memory[16'h3f83] <= 8'hb3;
		memory[16'h3f84] <= 8'he;
		memory[16'h3f85] <= 8'h2f;
		memory[16'h3f86] <= 8'hd2;
		memory[16'h3f87] <= 8'h17;
		memory[16'h3f88] <= 8'h29;
		memory[16'h3f89] <= 8'h9;
		memory[16'h3f8a] <= 8'h32;
		memory[16'h3f8b] <= 8'h12;
		memory[16'h3f8c] <= 8'h0;
		memory[16'h3f8d] <= 8'h6d;
		memory[16'h3f8e] <= 8'he6;
		memory[16'h3f8f] <= 8'h46;
		memory[16'h3f90] <= 8'h61;
		memory[16'h3f91] <= 8'hc3;
		memory[16'h3f92] <= 8'ha;
		memory[16'h3f93] <= 8'h7f;
		memory[16'h3f94] <= 8'h99;
		memory[16'h3f95] <= 8'hab;
		memory[16'h3f96] <= 8'he1;
		memory[16'h3f97] <= 8'h54;
		memory[16'h3f98] <= 8'h5d;
		memory[16'h3f99] <= 8'h63;
		memory[16'h3f9a] <= 8'h88;
		memory[16'h3f9b] <= 8'h86;
		memory[16'h3f9c] <= 8'hfc;
		memory[16'h3f9d] <= 8'he7;
		memory[16'h3f9e] <= 8'h32;
		memory[16'h3f9f] <= 8'h56;
		memory[16'h3fa0] <= 8'hb6;
		memory[16'h3fa1] <= 8'h4d;
		memory[16'h3fa2] <= 8'h9;
		memory[16'h3fa3] <= 8'hc4;
		memory[16'h3fa4] <= 8'h7d;
		memory[16'h3fa5] <= 8'hdb;
		memory[16'h3fa6] <= 8'hdc;
		memory[16'h3fa7] <= 8'ha6;
		memory[16'h3fa8] <= 8'he4;
		memory[16'h3fa9] <= 8'he;
		memory[16'h3faa] <= 8'hb8;
		memory[16'h3fab] <= 8'he4;
		memory[16'h3fac] <= 8'h7b;
		memory[16'h3fad] <= 8'h9e;
		memory[16'h3fae] <= 8'h2a;
		memory[16'h3faf] <= 8'hdd;
		memory[16'h3fb0] <= 8'h62;
		memory[16'h3fb1] <= 8'h34;
		memory[16'h3fb2] <= 8'h5c;
		memory[16'h3fb3] <= 8'hfb;
		memory[16'h3fb4] <= 8'hdf;
		memory[16'h3fb5] <= 8'h3e;
		memory[16'h3fb6] <= 8'h4f;
		memory[16'h3fb7] <= 8'h3d;
		memory[16'h3fb8] <= 8'ha1;
		memory[16'h3fb9] <= 8'hd8;
		memory[16'h3fba] <= 8'hc3;
		memory[16'h3fbb] <= 8'h9d;
		memory[16'h3fbc] <= 8'hbf;
		memory[16'h3fbd] <= 8'hf5;
		memory[16'h3fbe] <= 8'hf3;
		memory[16'h3fbf] <= 8'h75;
		memory[16'h3fc0] <= 8'h43;
		memory[16'h3fc1] <= 8'hfc;
		memory[16'h3fc2] <= 8'h3a;
		memory[16'h3fc3] <= 8'hc0;
		memory[16'h3fc4] <= 8'hd7;
		memory[16'h3fc5] <= 8'h16;
		memory[16'h3fc6] <= 8'h66;
		memory[16'h3fc7] <= 8'hbb;
		memory[16'h3fc8] <= 8'h24;
		memory[16'h3fc9] <= 8'h1e;
		memory[16'h3fca] <= 8'h9f;
		memory[16'h3fcb] <= 8'ha0;
		memory[16'h3fcc] <= 8'hbd;
		memory[16'h3fcd] <= 8'hca;
		memory[16'h3fce] <= 8'h7d;
		memory[16'h3fcf] <= 8'h1f;
		memory[16'h3fd0] <= 8'hfe;
		memory[16'h3fd1] <= 8'hd9;
		memory[16'h3fd2] <= 8'h1a;
		memory[16'h3fd3] <= 8'hde;
		memory[16'h3fd4] <= 8'h17;
		memory[16'h3fd5] <= 8'h6a;
		memory[16'h3fd6] <= 8'h1b;
		memory[16'h3fd7] <= 8'hb8;
		memory[16'h3fd8] <= 8'h42;
		memory[16'h3fd9] <= 8'hde;
		memory[16'h3fda] <= 8'h55;
		memory[16'h3fdb] <= 8'h1;
		memory[16'h3fdc] <= 8'hd4;
		memory[16'h3fdd] <= 8'h48;
		memory[16'h3fde] <= 8'h77;
		memory[16'h3fdf] <= 8'h17;
		memory[16'h3fe0] <= 8'h44;
		memory[16'h3fe1] <= 8'hb1;
		memory[16'h3fe2] <= 8'hd7;
		memory[16'h3fe3] <= 8'h1b;
		memory[16'h3fe4] <= 8'hc7;
		memory[16'h3fe5] <= 8'h3d;
		memory[16'h3fe6] <= 8'hd6;
		memory[16'h3fe7] <= 8'heb;
		memory[16'h3fe8] <= 8'h5b;
		memory[16'h3fe9] <= 8'h76;
		memory[16'h3fea] <= 8'h8b;
		memory[16'h3feb] <= 8'h18;
		memory[16'h3fec] <= 8'h40;
		memory[16'h3fed] <= 8'h8;
		memory[16'h3fee] <= 8'h37;
		memory[16'h3fef] <= 8'h3e;
		memory[16'h3ff0] <= 8'he2;
		memory[16'h3ff1] <= 8'h52;
		memory[16'h3ff2] <= 8'h1c;
		memory[16'h3ff3] <= 8'hf9;
		memory[16'h3ff4] <= 8'hbc;
		memory[16'h3ff5] <= 8'h37;
		memory[16'h3ff6] <= 8'hb2;
		memory[16'h3ff7] <= 8'hfe;
		memory[16'h3ff8] <= 8'h16;
		memory[16'h3ff9] <= 8'h7;
		memory[16'h3ffa] <= 8'hff;
		memory[16'h3ffb] <= 8'hea;
		memory[16'h3ffc] <= 8'h50;
		memory[16'h3ffd] <= 8'h76;
		memory[16'h3ffe] <= 8'h1;
		memory[16'h3fff] <= 8'h94;
		memory[16'h4000] <= 8'h27;
		memory[16'h4001] <= 8'hd8;
		memory[16'h4002] <= 8'hb0;
		memory[16'h4003] <= 8'hee;
		memory[16'h4004] <= 8'h15;
		memory[16'h4005] <= 8'h86;
		memory[16'h4006] <= 8'hda;
		memory[16'h4007] <= 8'h70;
		memory[16'h4008] <= 8'hfc;
		memory[16'h4009] <= 8'h65;
		memory[16'h400a] <= 8'h89;
		memory[16'h400b] <= 8'h3c;
		memory[16'h400c] <= 8'h6e;
		memory[16'h400d] <= 8'hc0;
		memory[16'h400e] <= 8'h7b;
		memory[16'h400f] <= 8'h50;
		memory[16'h4010] <= 8'h12;
		memory[16'h4011] <= 8'h97;
		memory[16'h4012] <= 8'h49;
		memory[16'h4013] <= 8'hce;
		memory[16'h4014] <= 8'hcf;
		memory[16'h4015] <= 8'hfb;
		memory[16'h4016] <= 8'hcc;
		memory[16'h4017] <= 8'he5;
		memory[16'h4018] <= 8'h3;
		memory[16'h4019] <= 8'hcc;
		memory[16'h401a] <= 8'hcf;
		memory[16'h401b] <= 8'h53;
		memory[16'h401c] <= 8'h42;
		memory[16'h401d] <= 8'hd0;
		memory[16'h401e] <= 8'he7;
		memory[16'h401f] <= 8'h6a;
		memory[16'h4020] <= 8'ha8;
		memory[16'h4021] <= 8'h97;
		memory[16'h4022] <= 8'h58;
		memory[16'h4023] <= 8'hbd;
		memory[16'h4024] <= 8'h1e;
		memory[16'h4025] <= 8'h32;
		memory[16'h4026] <= 8'h2d;
		memory[16'h4027] <= 8'h1a;
		memory[16'h4028] <= 8'h98;
		memory[16'h4029] <= 8'hb6;
		memory[16'h402a] <= 8'h57;
		memory[16'h402b] <= 8'h6;
		memory[16'h402c] <= 8'h77;
		memory[16'h402d] <= 8'hd2;
		memory[16'h402e] <= 8'h56;
		memory[16'h402f] <= 8'h89;
		memory[16'h4030] <= 8'h69;
		memory[16'h4031] <= 8'h9f;
		memory[16'h4032] <= 8'h58;
		memory[16'h4033] <= 8'h38;
		memory[16'h4034] <= 8'h9b;
		memory[16'h4035] <= 8'h24;
		memory[16'h4036] <= 8'h1d;
		memory[16'h4037] <= 8'h9e;
		memory[16'h4038] <= 8'hf0;
		memory[16'h4039] <= 8'hec;
		memory[16'h403a] <= 8'hf1;
		memory[16'h403b] <= 8'h33;
		memory[16'h403c] <= 8'hbc;
		memory[16'h403d] <= 8'hd8;
		memory[16'h403e] <= 8'h9d;
		memory[16'h403f] <= 8'h64;
		memory[16'h4040] <= 8'h70;
		memory[16'h4041] <= 8'hf5;
		memory[16'h4042] <= 8'h21;
		memory[16'h4043] <= 8'h8e;
		memory[16'h4044] <= 8'h28;
		memory[16'h4045] <= 8'h4f;
		memory[16'h4046] <= 8'ha8;
		memory[16'h4047] <= 8'hc0;
		memory[16'h4048] <= 8'h5;
		memory[16'h4049] <= 8'hff;
		memory[16'h404a] <= 8'hc6;
		memory[16'h404b] <= 8'h7c;
		memory[16'h404c] <= 8'hd1;
		memory[16'h404d] <= 8'h1c;
		memory[16'h404e] <= 8'h6;
		memory[16'h404f] <= 8'h3b;
		memory[16'h4050] <= 8'hbb;
		memory[16'h4051] <= 8'h5e;
		memory[16'h4052] <= 8'h73;
		memory[16'h4053] <= 8'h56;
		memory[16'h4054] <= 8'h82;
		memory[16'h4055] <= 8'h91;
		memory[16'h4056] <= 8'hf4;
		memory[16'h4057] <= 8'h73;
		memory[16'h4058] <= 8'h7d;
		memory[16'h4059] <= 8'he5;
		memory[16'h405a] <= 8'ha6;
		memory[16'h405b] <= 8'h3a;
		memory[16'h405c] <= 8'hbe;
		memory[16'h405d] <= 8'h43;
		memory[16'h405e] <= 8'h9e;
		memory[16'h405f] <= 8'h2e;
		memory[16'h4060] <= 8'h38;
		memory[16'h4061] <= 8'hc0;
		memory[16'h4062] <= 8'hbc;
		memory[16'h4063] <= 8'h60;
		memory[16'h4064] <= 8'hf;
		memory[16'h4065] <= 8'h64;
		memory[16'h4066] <= 8'h20;
		memory[16'h4067] <= 8'h14;
		memory[16'h4068] <= 8'h64;
		memory[16'h4069] <= 8'he6;
		memory[16'h406a] <= 8'h91;
		memory[16'h406b] <= 8'h35;
		memory[16'h406c] <= 8'h2;
		memory[16'h406d] <= 8'h97;
		memory[16'h406e] <= 8'h70;
		memory[16'h406f] <= 8'hbe;
		memory[16'h4070] <= 8'hf5;
		memory[16'h4071] <= 8'he4;
		memory[16'h4072] <= 8'h14;
		memory[16'h4073] <= 8'h77;
		memory[16'h4074] <= 8'h75;
		memory[16'h4075] <= 8'h9;
		memory[16'h4076] <= 8'hea;
		memory[16'h4077] <= 8'hf2;
		memory[16'h4078] <= 8'hee;
		memory[16'h4079] <= 8'h90;
		memory[16'h407a] <= 8'h2c;
		memory[16'h407b] <= 8'hac;
		memory[16'h407c] <= 8'hd3;
		memory[16'h407d] <= 8'hcb;
		memory[16'h407e] <= 8'hda;
		memory[16'h407f] <= 8'hc;
		memory[16'h4080] <= 8'h8b;
		memory[16'h4081] <= 8'h96;
		memory[16'h4082] <= 8'h6c;
		memory[16'h4083] <= 8'h9a;
		memory[16'h4084] <= 8'hfb;
		memory[16'h4085] <= 8'h8d;
		memory[16'h4086] <= 8'hae;
		memory[16'h4087] <= 8'h5f;
		memory[16'h4088] <= 8'h73;
		memory[16'h4089] <= 8'h3f;
		memory[16'h408a] <= 8'h94;
		memory[16'h408b] <= 8'h76;
		memory[16'h408c] <= 8'hd6;
		memory[16'h408d] <= 8'h5;
		memory[16'h408e] <= 8'h34;
		memory[16'h408f] <= 8'hcb;
		memory[16'h4090] <= 8'he9;
		memory[16'h4091] <= 8'h48;
		memory[16'h4092] <= 8'h43;
		memory[16'h4093] <= 8'h5e;
		memory[16'h4094] <= 8'h51;
		memory[16'h4095] <= 8'h2d;
		memory[16'h4096] <= 8'h50;
		memory[16'h4097] <= 8'h40;
		memory[16'h4098] <= 8'hbe;
		memory[16'h4099] <= 8'h7d;
		memory[16'h409a] <= 8'hec;
		memory[16'h409b] <= 8'h91;
		memory[16'h409c] <= 8'h48;
		memory[16'h409d] <= 8'hc7;
		memory[16'h409e] <= 8'h9d;
		memory[16'h409f] <= 8'hd3;
		memory[16'h40a0] <= 8'h5d;
		memory[16'h40a1] <= 8'ha;
		memory[16'h40a2] <= 8'h6d;
		memory[16'h40a3] <= 8'h58;
		memory[16'h40a4] <= 8'h97;
		memory[16'h40a5] <= 8'h1b;
		memory[16'h40a6] <= 8'hb7;
		memory[16'h40a7] <= 8'ha;
		memory[16'h40a8] <= 8'h5b;
		memory[16'h40a9] <= 8'h4c;
		memory[16'h40aa] <= 8'h80;
		memory[16'h40ab] <= 8'h31;
		memory[16'h40ac] <= 8'h51;
		memory[16'h40ad] <= 8'hb4;
		memory[16'h40ae] <= 8'hfd;
		memory[16'h40af] <= 8'h3a;
		memory[16'h40b0] <= 8'hfd;
		memory[16'h40b1] <= 8'h40;
		memory[16'h40b2] <= 8'h98;
		memory[16'h40b3] <= 8'h4e;
		memory[16'h40b4] <= 8'h6d;
		memory[16'h40b5] <= 8'he8;
		memory[16'h40b6] <= 8'h8e;
		memory[16'h40b7] <= 8'h2b;
		memory[16'h40b8] <= 8'h65;
		memory[16'h40b9] <= 8'h7b;
		memory[16'h40ba] <= 8'hbd;
		memory[16'h40bb] <= 8'had;
		memory[16'h40bc] <= 8'h42;
		memory[16'h40bd] <= 8'h5a;
		memory[16'h40be] <= 8'h80;
		memory[16'h40bf] <= 8'h9f;
		memory[16'h40c0] <= 8'h64;
		memory[16'h40c1] <= 8'hed;
		memory[16'h40c2] <= 8'hf8;
		memory[16'h40c3] <= 8'hfb;
		memory[16'h40c4] <= 8'h9;
		memory[16'h40c5] <= 8'haf;
		memory[16'h40c6] <= 8'h6;
		memory[16'h40c7] <= 8'h64;
		memory[16'h40c8] <= 8'hfb;
		memory[16'h40c9] <= 8'h86;
		memory[16'h40ca] <= 8'h95;
		memory[16'h40cb] <= 8'h4c;
		memory[16'h40cc] <= 8'h3b;
		memory[16'h40cd] <= 8'h92;
		memory[16'h40ce] <= 8'h86;
		memory[16'h40cf] <= 8'h38;
		memory[16'h40d0] <= 8'hd2;
		memory[16'h40d1] <= 8'h1e;
		memory[16'h40d2] <= 8'h86;
		memory[16'h40d3] <= 8'h40;
		memory[16'h40d4] <= 8'h7;
		memory[16'h40d5] <= 8'h15;
		memory[16'h40d6] <= 8'h6b;
		memory[16'h40d7] <= 8'h6c;
		memory[16'h40d8] <= 8'h90;
		memory[16'h40d9] <= 8'h28;
		memory[16'h40da] <= 8'h1a;
		memory[16'h40db] <= 8'hd2;
		memory[16'h40dc] <= 8'h83;
		memory[16'h40dd] <= 8'h9a;
		memory[16'h40de] <= 8'h71;
		memory[16'h40df] <= 8'he7;
		memory[16'h40e0] <= 8'h88;
		memory[16'h40e1] <= 8'h69;
		memory[16'h40e2] <= 8'he3;
		memory[16'h40e3] <= 8'h91;
		memory[16'h40e4] <= 8'h19;
		memory[16'h40e5] <= 8'he9;
		memory[16'h40e6] <= 8'hf5;
		memory[16'h40e7] <= 8'h14;
		memory[16'h40e8] <= 8'h6f;
		memory[16'h40e9] <= 8'h8a;
		memory[16'h40ea] <= 8'h61;
		memory[16'h40eb] <= 8'haa;
		memory[16'h40ec] <= 8'h1d;
		memory[16'h40ed] <= 8'he7;
		memory[16'h40ee] <= 8'he2;
		memory[16'h40ef] <= 8'hef;
		memory[16'h40f0] <= 8'h6;
		memory[16'h40f1] <= 8'h69;
		memory[16'h40f2] <= 8'h2f;
		memory[16'h40f3] <= 8'hd;
		memory[16'h40f4] <= 8'h7e;
		memory[16'h40f5] <= 8'h9b;
		memory[16'h40f6] <= 8'h79;
		memory[16'h40f7] <= 8'he;
		memory[16'h40f8] <= 8'hc3;
		memory[16'h40f9] <= 8'h93;
		memory[16'h40fa] <= 8'he0;
		memory[16'h40fb] <= 8'h46;
		memory[16'h40fc] <= 8'h2e;
		memory[16'h40fd] <= 8'h51;
		memory[16'h40fe] <= 8'h2e;
		memory[16'h40ff] <= 8'hb6;
		memory[16'h4100] <= 8'hbb;
		memory[16'h4101] <= 8'h11;
		memory[16'h4102] <= 8'h47;
		memory[16'h4103] <= 8'hd4;
		memory[16'h4104] <= 8'hfa;
		memory[16'h4105] <= 8'h3c;
		memory[16'h4106] <= 8'he8;
		memory[16'h4107] <= 8'h69;
		memory[16'h4108] <= 8'hc6;
		memory[16'h4109] <= 8'h49;
		memory[16'h410a] <= 8'h14;
		memory[16'h410b] <= 8'he3;
		memory[16'h410c] <= 8'h31;
		memory[16'h410d] <= 8'hf6;
		memory[16'h410e] <= 8'hd3;
		memory[16'h410f] <= 8'h37;
		memory[16'h4110] <= 8'h5f;
		memory[16'h4111] <= 8'h2;
		memory[16'h4112] <= 8'h44;
		memory[16'h4113] <= 8'hdd;
		memory[16'h4114] <= 8'h9d;
		memory[16'h4115] <= 8'hbd;
		memory[16'h4116] <= 8'heb;
		memory[16'h4117] <= 8'h61;
		memory[16'h4118] <= 8'h51;
		memory[16'h4119] <= 8'hcb;
		memory[16'h411a] <= 8'ha7;
		memory[16'h411b] <= 8'h7f;
		memory[16'h411c] <= 8'h1d;
		memory[16'h411d] <= 8'hd5;
		memory[16'h411e] <= 8'h35;
		memory[16'h411f] <= 8'hd8;
		memory[16'h4120] <= 8'he6;
		memory[16'h4121] <= 8'h7c;
		memory[16'h4122] <= 8'hac;
		memory[16'h4123] <= 8'he0;
		memory[16'h4124] <= 8'hb8;
		memory[16'h4125] <= 8'h94;
		memory[16'h4126] <= 8'h4a;
		memory[16'h4127] <= 8'h7e;
		memory[16'h4128] <= 8'hde;
		memory[16'h4129] <= 8'h5e;
		memory[16'h412a] <= 8'h62;
		memory[16'h412b] <= 8'hf;
		memory[16'h412c] <= 8'h54;
		memory[16'h412d] <= 8'h35;
		memory[16'h412e] <= 8'h46;
		memory[16'h412f] <= 8'hb4;
		memory[16'h4130] <= 8'h37;
		memory[16'h4131] <= 8'h8a;
		memory[16'h4132] <= 8'h91;
		memory[16'h4133] <= 8'hd5;
		memory[16'h4134] <= 8'h47;
		memory[16'h4135] <= 8'h7d;
		memory[16'h4136] <= 8'h36;
		memory[16'h4137] <= 8'h98;
		memory[16'h4138] <= 8'h48;
		memory[16'h4139] <= 8'hdd;
		memory[16'h413a] <= 8'h17;
		memory[16'h413b] <= 8'h65;
		memory[16'h413c] <= 8'hb3;
		memory[16'h413d] <= 8'h4c;
		memory[16'h413e] <= 8'h3d;
		memory[16'h413f] <= 8'h99;
		memory[16'h4140] <= 8'hc8;
		memory[16'h4141] <= 8'he9;
		memory[16'h4142] <= 8'h7a;
		memory[16'h4143] <= 8'h80;
		memory[16'h4144] <= 8'h7e;
		memory[16'h4145] <= 8'hc4;
		memory[16'h4146] <= 8'hff;
		memory[16'h4147] <= 8'h5c;
		memory[16'h4148] <= 8'h22;
		memory[16'h4149] <= 8'h61;
		memory[16'h414a] <= 8'h6b;
		memory[16'h414b] <= 8'h76;
		memory[16'h414c] <= 8'h96;
		memory[16'h414d] <= 8'hb1;
		memory[16'h414e] <= 8'h2a;
		memory[16'h414f] <= 8'hcd;
		memory[16'h4150] <= 8'h3b;
		memory[16'h4151] <= 8'hbc;
		memory[16'h4152] <= 8'ha2;
		memory[16'h4153] <= 8'h82;
		memory[16'h4154] <= 8'h39;
		memory[16'h4155] <= 8'hd8;
		memory[16'h4156] <= 8'h1b;
		memory[16'h4157] <= 8'h81;
		memory[16'h4158] <= 8'hb6;
		memory[16'h4159] <= 8'h32;
		memory[16'h415a] <= 8'he7;
		memory[16'h415b] <= 8'h69;
		memory[16'h415c] <= 8'h7f;
		memory[16'h415d] <= 8'h24;
		memory[16'h415e] <= 8'h2;
		memory[16'h415f] <= 8'h47;
		memory[16'h4160] <= 8'he;
		memory[16'h4161] <= 8'h7c;
		memory[16'h4162] <= 8'hc8;
		memory[16'h4163] <= 8'h8c;
		memory[16'h4164] <= 8'h40;
		memory[16'h4165] <= 8'hc7;
		memory[16'h4166] <= 8'he8;
		memory[16'h4167] <= 8'h62;
		memory[16'h4168] <= 8'h28;
		memory[16'h4169] <= 8'h53;
		memory[16'h416a] <= 8'hd9;
		memory[16'h416b] <= 8'hbe;
		memory[16'h416c] <= 8'h4;
		memory[16'h416d] <= 8'h3;
		memory[16'h416e] <= 8'h8b;
		memory[16'h416f] <= 8'h3f;
		memory[16'h4170] <= 8'hbf;
		memory[16'h4171] <= 8'h2e;
		memory[16'h4172] <= 8'hc1;
		memory[16'h4173] <= 8'hf8;
		memory[16'h4174] <= 8'h6;
		memory[16'h4175] <= 8'hdc;
		memory[16'h4176] <= 8'h7a;
		memory[16'h4177] <= 8'hbc;
		memory[16'h4178] <= 8'hf;
		memory[16'h4179] <= 8'h61;
		memory[16'h417a] <= 8'h25;
		memory[16'h417b] <= 8'h8e;
		memory[16'h417c] <= 8'h85;
		memory[16'h417d] <= 8'h28;
		memory[16'h417e] <= 8'hd5;
		memory[16'h417f] <= 8'h93;
		memory[16'h4180] <= 8'ha4;
		memory[16'h4181] <= 8'h9d;
		memory[16'h4182] <= 8'h1f;
		memory[16'h4183] <= 8'he5;
		memory[16'h4184] <= 8'h64;
		memory[16'h4185] <= 8'h7;
		memory[16'h4186] <= 8'h47;
		memory[16'h4187] <= 8'h8c;
		memory[16'h4188] <= 8'h5a;
		memory[16'h4189] <= 8'h20;
		memory[16'h418a] <= 8'h4a;
		memory[16'h418b] <= 8'h5e;
		memory[16'h418c] <= 8'h24;
		memory[16'h418d] <= 8'hd6;
		memory[16'h418e] <= 8'h9d;
		memory[16'h418f] <= 8'he3;
		memory[16'h4190] <= 8'h4;
		memory[16'h4191] <= 8'h5f;
		memory[16'h4192] <= 8'hdc;
		memory[16'h4193] <= 8'ha;
		memory[16'h4194] <= 8'h3b;
		memory[16'h4195] <= 8'h56;
		memory[16'h4196] <= 8'hc7;
		memory[16'h4197] <= 8'h4a;
		memory[16'h4198] <= 8'hb7;
		memory[16'h4199] <= 8'hec;
		memory[16'h419a] <= 8'hd8;
		memory[16'h419b] <= 8'h3c;
		memory[16'h419c] <= 8'h14;
		memory[16'h419d] <= 8'hae;
		memory[16'h419e] <= 8'hd0;
		memory[16'h419f] <= 8'hb9;
		memory[16'h41a0] <= 8'h4b;
		memory[16'h41a1] <= 8'hef;
		memory[16'h41a2] <= 8'h9e;
		memory[16'h41a3] <= 8'hb0;
		memory[16'h41a4] <= 8'hf7;
		memory[16'h41a5] <= 8'he5;
		memory[16'h41a6] <= 8'h3c;
		memory[16'h41a7] <= 8'h51;
		memory[16'h41a8] <= 8'h6;
		memory[16'h41a9] <= 8'h87;
		memory[16'h41aa] <= 8'hb0;
		memory[16'h41ab] <= 8'h2a;
		memory[16'h41ac] <= 8'h5d;
		memory[16'h41ad] <= 8'h4d;
		memory[16'h41ae] <= 8'hd;
		memory[16'h41af] <= 8'h61;
		memory[16'h41b0] <= 8'hac;
		memory[16'h41b1] <= 8'he9;
		memory[16'h41b2] <= 8'h6b;
		memory[16'h41b3] <= 8'he8;
		memory[16'h41b4] <= 8'h3f;
		memory[16'h41b5] <= 8'h32;
		memory[16'h41b6] <= 8'h32;
		memory[16'h41b7] <= 8'hf6;
		memory[16'h41b8] <= 8'h1f;
		memory[16'h41b9] <= 8'hb;
		memory[16'h41ba] <= 8'h33;
		memory[16'h41bb] <= 8'h33;
		memory[16'h41bc] <= 8'hb9;
		memory[16'h41bd] <= 8'h3;
		memory[16'h41be] <= 8'hec;
		memory[16'h41bf] <= 8'h4;
		memory[16'h41c0] <= 8'hf2;
		memory[16'h41c1] <= 8'h8a;
		memory[16'h41c2] <= 8'hb4;
		memory[16'h41c3] <= 8'he9;
		memory[16'h41c4] <= 8'h70;
		memory[16'h41c5] <= 8'hf1;
		memory[16'h41c6] <= 8'h3b;
		memory[16'h41c7] <= 8'h76;
		memory[16'h41c8] <= 8'h78;
		memory[16'h41c9] <= 8'heb;
		memory[16'h41ca] <= 8'ha0;
		memory[16'h41cb] <= 8'hd5;
		memory[16'h41cc] <= 8'h38;
		memory[16'h41cd] <= 8'had;
		memory[16'h41ce] <= 8'h36;
		memory[16'h41cf] <= 8'he5;
		memory[16'h41d0] <= 8'h97;
		memory[16'h41d1] <= 8'ha1;
		memory[16'h41d2] <= 8'hcd;
		memory[16'h41d3] <= 8'hd6;
		memory[16'h41d4] <= 8'hd4;
		memory[16'h41d5] <= 8'hff;
		memory[16'h41d6] <= 8'hcd;
		memory[16'h41d7] <= 8'hf3;
		memory[16'h41d8] <= 8'ha;
		memory[16'h41d9] <= 8'h0;
		memory[16'h41da] <= 8'h26;
		memory[16'h41db] <= 8'hc3;
		memory[16'h41dc] <= 8'h3;
		memory[16'h41dd] <= 8'h13;
		memory[16'h41de] <= 8'hc8;
		memory[16'h41df] <= 8'hf5;
		memory[16'h41e0] <= 8'h9d;
		memory[16'h41e1] <= 8'h7c;
		memory[16'h41e2] <= 8'hdf;
		memory[16'h41e3] <= 8'hd;
		memory[16'h41e4] <= 8'h6d;
		memory[16'h41e5] <= 8'h1a;
		memory[16'h41e6] <= 8'h83;
		memory[16'h41e7] <= 8'he5;
		memory[16'h41e8] <= 8'h5;
		memory[16'h41e9] <= 8'h23;
		memory[16'h41ea] <= 8'hba;
		memory[16'h41eb] <= 8'h3d;
		memory[16'h41ec] <= 8'hd1;
		memory[16'h41ed] <= 8'hf0;
		memory[16'h41ee] <= 8'h22;
		memory[16'h41ef] <= 8'h68;
		memory[16'h41f0] <= 8'h92;
		memory[16'h41f1] <= 8'hef;
		memory[16'h41f2] <= 8'h3e;
		memory[16'h41f3] <= 8'h66;
		memory[16'h41f4] <= 8'hef;
		memory[16'h41f5] <= 8'hb;
		memory[16'h41f6] <= 8'h59;
		memory[16'h41f7] <= 8'hf9;
		memory[16'h41f8] <= 8'hb;
		memory[16'h41f9] <= 8'h7f;
		memory[16'h41fa] <= 8'hbd;
		memory[16'h41fb] <= 8'he;
		memory[16'h41fc] <= 8'h92;
		memory[16'h41fd] <= 8'h85;
		memory[16'h41fe] <= 8'h4;
		memory[16'h41ff] <= 8'h30;
		memory[16'h4200] <= 8'h1;
		memory[16'h4201] <= 8'he3;
		memory[16'h4202] <= 8'h3d;
		memory[16'h4203] <= 8'h6f;
		memory[16'h4204] <= 8'hfd;
		memory[16'h4205] <= 8'hc1;
		memory[16'h4206] <= 8'h54;
		memory[16'h4207] <= 8'h2;
		memory[16'h4208] <= 8'he4;
		memory[16'h4209] <= 8'hf;
		memory[16'h420a] <= 8'h3f;
		memory[16'h420b] <= 8'hb5;
		memory[16'h420c] <= 8'hff;
		memory[16'h420d] <= 8'h62;
		memory[16'h420e] <= 8'h1d;
		memory[16'h420f] <= 8'h91;
		memory[16'h4210] <= 8'h51;
		memory[16'h4211] <= 8'h5c;
		memory[16'h4212] <= 8'hf7;
		memory[16'h4213] <= 8'h40;
		memory[16'h4214] <= 8'h67;
		memory[16'h4215] <= 8'h50;
		memory[16'h4216] <= 8'h3a;
		memory[16'h4217] <= 8'h73;
		memory[16'h4218] <= 8'hd0;
		memory[16'h4219] <= 8'hf7;
		memory[16'h421a] <= 8'h81;
		memory[16'h421b] <= 8'h62;
		memory[16'h421c] <= 8'h7c;
		memory[16'h421d] <= 8'h85;
		memory[16'h421e] <= 8'h92;
		memory[16'h421f] <= 8'h7d;
		memory[16'h4220] <= 8'h68;
		memory[16'h4221] <= 8'hd0;
		memory[16'h4222] <= 8'hec;
		memory[16'h4223] <= 8'h65;
		memory[16'h4224] <= 8'h91;
		memory[16'h4225] <= 8'h41;
		memory[16'h4226] <= 8'h67;
		memory[16'h4227] <= 8'h75;
		memory[16'h4228] <= 8'h50;
		memory[16'h4229] <= 8'ha7;
		memory[16'h422a] <= 8'h2b;
		memory[16'h422b] <= 8'h4f;
		memory[16'h422c] <= 8'h9;
		memory[16'h422d] <= 8'h48;
		memory[16'h422e] <= 8'he1;
		memory[16'h422f] <= 8'h5a;
		memory[16'h4230] <= 8'ha4;
		memory[16'h4231] <= 8'hd8;
		memory[16'h4232] <= 8'h9b;
		memory[16'h4233] <= 8'hc;
		memory[16'h4234] <= 8'h29;
		memory[16'h4235] <= 8'hd5;
		memory[16'h4236] <= 8'h7f;
		memory[16'h4237] <= 8'hf9;
		memory[16'h4238] <= 8'hcc;
		memory[16'h4239] <= 8'h0;
		memory[16'h423a] <= 8'h5b;
		memory[16'h423b] <= 8'h48;
		memory[16'h423c] <= 8'h86;
		memory[16'h423d] <= 8'hee;
		memory[16'h423e] <= 8'hc5;
		memory[16'h423f] <= 8'hee;
		memory[16'h4240] <= 8'hbe;
		memory[16'h4241] <= 8'hb2;
		memory[16'h4242] <= 8'h54;
		memory[16'h4243] <= 8'h4f;
		memory[16'h4244] <= 8'hf3;
		memory[16'h4245] <= 8'hbb;
		memory[16'h4246] <= 8'hc4;
		memory[16'h4247] <= 8'h43;
		memory[16'h4248] <= 8'h62;
		memory[16'h4249] <= 8'hef;
		memory[16'h424a] <= 8'h92;
		memory[16'h424b] <= 8'h6b;
		memory[16'h424c] <= 8'h38;
		memory[16'h424d] <= 8'h73;
		memory[16'h424e] <= 8'hc6;
		memory[16'h424f] <= 8'hdc;
		memory[16'h4250] <= 8'h4c;
		memory[16'h4251] <= 8'h61;
		memory[16'h4252] <= 8'he8;
		memory[16'h4253] <= 8'h75;
		memory[16'h4254] <= 8'h36;
		memory[16'h4255] <= 8'h67;
		memory[16'h4256] <= 8'h6e;
		memory[16'h4257] <= 8'h2;
		memory[16'h4258] <= 8'h68;
		memory[16'h4259] <= 8'hc9;
		memory[16'h425a] <= 8'h4a;
		memory[16'h425b] <= 8'hee;
		memory[16'h425c] <= 8'hb7;
		memory[16'h425d] <= 8'hf;
		memory[16'h425e] <= 8'hdc;
		memory[16'h425f] <= 8'h75;
		memory[16'h4260] <= 8'hc1;
		memory[16'h4261] <= 8'h30;
		memory[16'h4262] <= 8'hc4;
		memory[16'h4263] <= 8'hb4;
		memory[16'h4264] <= 8'hec;
		memory[16'h4265] <= 8'h89;
		memory[16'h4266] <= 8'hf7;
		memory[16'h4267] <= 8'h4e;
		memory[16'h4268] <= 8'h78;
		memory[16'h4269] <= 8'h8a;
		memory[16'h426a] <= 8'hba;
		memory[16'h426b] <= 8'hb0;
		memory[16'h426c] <= 8'hfd;
		memory[16'h426d] <= 8'h80;
		memory[16'h426e] <= 8'h8d;
		memory[16'h426f] <= 8'h49;
		memory[16'h4270] <= 8'he1;
		memory[16'h4271] <= 8'h75;
		memory[16'h4272] <= 8'hbe;
		memory[16'h4273] <= 8'h17;
		memory[16'h4274] <= 8'hdd;
		memory[16'h4275] <= 8'h2c;
		memory[16'h4276] <= 8'h19;
		memory[16'h4277] <= 8'h45;
		memory[16'h4278] <= 8'hf6;
		memory[16'h4279] <= 8'h63;
		memory[16'h427a] <= 8'h33;
		memory[16'h427b] <= 8'had;
		memory[16'h427c] <= 8'h72;
		memory[16'h427d] <= 8'hf;
		memory[16'h427e] <= 8'h23;
		memory[16'h427f] <= 8'h34;
		memory[16'h4280] <= 8'h40;
		memory[16'h4281] <= 8'he7;
		memory[16'h4282] <= 8'he8;
		memory[16'h4283] <= 8'h2c;
		memory[16'h4284] <= 8'h70;
		memory[16'h4285] <= 8'he0;
		memory[16'h4286] <= 8'h7a;
		memory[16'h4287] <= 8'he9;
		memory[16'h4288] <= 8'h6a;
		memory[16'h4289] <= 8'h34;
		memory[16'h428a] <= 8'h99;
		memory[16'h428b] <= 8'h67;
		memory[16'h428c] <= 8'hb4;
		memory[16'h428d] <= 8'h26;
		memory[16'h428e] <= 8'hb1;
		memory[16'h428f] <= 8'h95;
		memory[16'h4290] <= 8'h9c;
		memory[16'h4291] <= 8'h6f;
		memory[16'h4292] <= 8'hac;
		memory[16'h4293] <= 8'h79;
		memory[16'h4294] <= 8'h9c;
		memory[16'h4295] <= 8'hc5;
		memory[16'h4296] <= 8'hbe;
		memory[16'h4297] <= 8'h92;
		memory[16'h4298] <= 8'h28;
		memory[16'h4299] <= 8'hf1;
		memory[16'h429a] <= 8'h3f;
		memory[16'h429b] <= 8'h9b;
		memory[16'h429c] <= 8'h0;
		memory[16'h429d] <= 8'h62;
		memory[16'h429e] <= 8'hcf;
		memory[16'h429f] <= 8'h40;
		memory[16'h42a0] <= 8'h4a;
		memory[16'h42a1] <= 8'hb7;
		memory[16'h42a2] <= 8'h6c;
		memory[16'h42a3] <= 8'hba;
		memory[16'h42a4] <= 8'h97;
		memory[16'h42a5] <= 8'he7;
		memory[16'h42a6] <= 8'ha3;
		memory[16'h42a7] <= 8'h1;
		memory[16'h42a8] <= 8'h1b;
		memory[16'h42a9] <= 8'h3d;
		memory[16'h42aa] <= 8'h69;
		memory[16'h42ab] <= 8'hd0;
		memory[16'h42ac] <= 8'h63;
		memory[16'h42ad] <= 8'h1a;
		memory[16'h42ae] <= 8'h65;
		memory[16'h42af] <= 8'hff;
		memory[16'h42b0] <= 8'h89;
		memory[16'h42b1] <= 8'h12;
		memory[16'h42b2] <= 8'h78;
		memory[16'h42b3] <= 8'h25;
		memory[16'h42b4] <= 8'hd7;
		memory[16'h42b5] <= 8'h36;
		memory[16'h42b6] <= 8'hb7;
		memory[16'h42b7] <= 8'h0;
		memory[16'h42b8] <= 8'h27;
		memory[16'h42b9] <= 8'hf7;
		memory[16'h42ba] <= 8'h9b;
		memory[16'h42bb] <= 8'h28;
		memory[16'h42bc] <= 8'h59;
		memory[16'h42bd] <= 8'h6a;
		memory[16'h42be] <= 8'h68;
		memory[16'h42bf] <= 8'ha3;
		memory[16'h42c0] <= 8'h21;
		memory[16'h42c1] <= 8'hd5;
		memory[16'h42c2] <= 8'h5e;
		memory[16'h42c3] <= 8'hb9;
		memory[16'h42c4] <= 8'hbc;
		memory[16'h42c5] <= 8'h1;
		memory[16'h42c6] <= 8'hba;
		memory[16'h42c7] <= 8'hd7;
		memory[16'h42c8] <= 8'h3e;
		memory[16'h42c9] <= 8'h23;
		memory[16'h42ca] <= 8'ha7;
		memory[16'h42cb] <= 8'ha2;
		memory[16'h42cc] <= 8'h3d;
		memory[16'h42cd] <= 8'hd;
		memory[16'h42ce] <= 8'ha1;
		memory[16'h42cf] <= 8'hc7;
		memory[16'h42d0] <= 8'h1f;
		memory[16'h42d1] <= 8'h1a;
		memory[16'h42d2] <= 8'hec;
		memory[16'h42d3] <= 8'hf6;
		memory[16'h42d4] <= 8'h50;
		memory[16'h42d5] <= 8'ha4;
		memory[16'h42d6] <= 8'hf6;
		memory[16'h42d7] <= 8'h78;
		memory[16'h42d8] <= 8'h9b;
		memory[16'h42d9] <= 8'h91;
		memory[16'h42da] <= 8'ha0;
		memory[16'h42db] <= 8'hf4;
		memory[16'h42dc] <= 8'hfb;
		memory[16'h42dd] <= 8'h8;
		memory[16'h42de] <= 8'h98;
		memory[16'h42df] <= 8'h1d;
		memory[16'h42e0] <= 8'hdd;
		memory[16'h42e1] <= 8'hf6;
		memory[16'h42e2] <= 8'hd6;
		memory[16'h42e3] <= 8'h99;
		memory[16'h42e4] <= 8'hf7;
		memory[16'h42e5] <= 8'h90;
		memory[16'h42e6] <= 8'h71;
		memory[16'h42e7] <= 8'h36;
		memory[16'h42e8] <= 8'hb4;
		memory[16'h42e9] <= 8'h18;
		memory[16'h42ea] <= 8'hd8;
		memory[16'h42eb] <= 8'hf1;
		memory[16'h42ec] <= 8'h25;
		memory[16'h42ed] <= 8'h79;
		memory[16'h42ee] <= 8'hb8;
		memory[16'h42ef] <= 8'h44;
		memory[16'h42f0] <= 8'h93;
		memory[16'h42f1] <= 8'ha5;
		memory[16'h42f2] <= 8'h3b;
		memory[16'h42f3] <= 8'he4;
		memory[16'h42f4] <= 8'h49;
		memory[16'h42f5] <= 8'h31;
		memory[16'h42f6] <= 8'h5c;
		memory[16'h42f7] <= 8'he4;
		memory[16'h42f8] <= 8'hc3;
		memory[16'h42f9] <= 8'hfc;
		memory[16'h42fa] <= 8'hd8;
		memory[16'h42fb] <= 8'hbe;
		memory[16'h42fc] <= 8'h4;
		memory[16'h42fd] <= 8'h70;
		memory[16'h42fe] <= 8'hdb;
		memory[16'h42ff] <= 8'he2;
		memory[16'h4300] <= 8'h66;
		memory[16'h4301] <= 8'hb1;
		memory[16'h4302] <= 8'h7b;
		memory[16'h4303] <= 8'h5e;
		memory[16'h4304] <= 8'h42;
		memory[16'h4305] <= 8'hec;
		memory[16'h4306] <= 8'h94;
		memory[16'h4307] <= 8'hf6;
		memory[16'h4308] <= 8'h5;
		memory[16'h4309] <= 8'h6c;
		memory[16'h430a] <= 8'he7;
		memory[16'h430b] <= 8'h2a;
		memory[16'h430c] <= 8'he5;
		memory[16'h430d] <= 8'ha0;
		memory[16'h430e] <= 8'h6f;
		memory[16'h430f] <= 8'h79;
		memory[16'h4310] <= 8'h45;
		memory[16'h4311] <= 8'haa;
		memory[16'h4312] <= 8'h5d;
		memory[16'h4313] <= 8'h8e;
		memory[16'h4314] <= 8'hdb;
		memory[16'h4315] <= 8'hb9;
		memory[16'h4316] <= 8'h72;
		memory[16'h4317] <= 8'h9e;
		memory[16'h4318] <= 8'hb5;
		memory[16'h4319] <= 8'h4a;
		memory[16'h431a] <= 8'h5d;
		memory[16'h431b] <= 8'hb9;
		memory[16'h431c] <= 8'hbb;
		memory[16'h431d] <= 8'h38;
		memory[16'h431e] <= 8'h9b;
		memory[16'h431f] <= 8'h21;
		memory[16'h4320] <= 8'hea;
		memory[16'h4321] <= 8'h17;
		memory[16'h4322] <= 8'h7f;
		memory[16'h4323] <= 8'h2c;
		memory[16'h4324] <= 8'h3;
		memory[16'h4325] <= 8'h13;
		memory[16'h4326] <= 8'h22;
		memory[16'h4327] <= 8'h8;
		memory[16'h4328] <= 8'h7f;
		memory[16'h4329] <= 8'h9;
		memory[16'h432a] <= 8'h33;
		memory[16'h432b] <= 8'h65;
		memory[16'h432c] <= 8'ha9;
		memory[16'h432d] <= 8'ha2;
		memory[16'h432e] <= 8'hde;
		memory[16'h432f] <= 8'hee;
		memory[16'h4330] <= 8'h4c;
		memory[16'h4331] <= 8'h3b;
		memory[16'h4332] <= 8'h7c;
		memory[16'h4333] <= 8'h27;
		memory[16'h4334] <= 8'hf4;
		memory[16'h4335] <= 8'hee;
		memory[16'h4336] <= 8'hc6;
		memory[16'h4337] <= 8'ha9;
		memory[16'h4338] <= 8'h39;
		memory[16'h4339] <= 8'h23;
		memory[16'h433a] <= 8'h62;
		memory[16'h433b] <= 8'hf4;
		memory[16'h433c] <= 8'h5b;
		memory[16'h433d] <= 8'hfe;
		memory[16'h433e] <= 8'h15;
		memory[16'h433f] <= 8'h45;
		memory[16'h4340] <= 8'h15;
		memory[16'h4341] <= 8'h95;
		memory[16'h4342] <= 8'h71;
		memory[16'h4343] <= 8'h18;
		memory[16'h4344] <= 8'ha8;
		memory[16'h4345] <= 8'h93;
		memory[16'h4346] <= 8'h21;
		memory[16'h4347] <= 8'h28;
		memory[16'h4348] <= 8'h9d;
		memory[16'h4349] <= 8'h54;
		memory[16'h434a] <= 8'h8d;
		memory[16'h434b] <= 8'h46;
		memory[16'h434c] <= 8'hf6;
		memory[16'h434d] <= 8'h6b;
		memory[16'h434e] <= 8'h35;
		memory[16'h434f] <= 8'h42;
		memory[16'h4350] <= 8'ha6;
		memory[16'h4351] <= 8'hb1;
		memory[16'h4352] <= 8'h69;
		memory[16'h4353] <= 8'h9a;
		memory[16'h4354] <= 8'ha0;
		memory[16'h4355] <= 8'h2f;
		memory[16'h4356] <= 8'h43;
		memory[16'h4357] <= 8'hd9;
		memory[16'h4358] <= 8'h52;
		memory[16'h4359] <= 8'ha5;
		memory[16'h435a] <= 8'hcd;
		memory[16'h435b] <= 8'hae;
		memory[16'h435c] <= 8'ha3;
		memory[16'h435d] <= 8'he2;
		memory[16'h435e] <= 8'hf3;
		memory[16'h435f] <= 8'hb8;
		memory[16'h4360] <= 8'h77;
		memory[16'h4361] <= 8'h65;
		memory[16'h4362] <= 8'hd1;
		memory[16'h4363] <= 8'h20;
		memory[16'h4364] <= 8'hf8;
		memory[16'h4365] <= 8'hf2;
		memory[16'h4366] <= 8'h48;
		memory[16'h4367] <= 8'h95;
		memory[16'h4368] <= 8'h46;
		memory[16'h4369] <= 8'hd5;
		memory[16'h436a] <= 8'hdc;
		memory[16'h436b] <= 8'h3c;
		memory[16'h436c] <= 8'h40;
		memory[16'h436d] <= 8'h11;
		memory[16'h436e] <= 8'h7e;
		memory[16'h436f] <= 8'he6;
		memory[16'h4370] <= 8'hc2;
		memory[16'h4371] <= 8'he7;
		memory[16'h4372] <= 8'h80;
		memory[16'h4373] <= 8'h62;
		memory[16'h4374] <= 8'h17;
		memory[16'h4375] <= 8'hc3;
		memory[16'h4376] <= 8'h3b;
		memory[16'h4377] <= 8'h69;
		memory[16'h4378] <= 8'h68;
		memory[16'h4379] <= 8'h8;
		memory[16'h437a] <= 8'h17;
		memory[16'h437b] <= 8'hc;
		memory[16'h437c] <= 8'heb;
		memory[16'h437d] <= 8'hb;
		memory[16'h437e] <= 8'hc4;
		memory[16'h437f] <= 8'h62;
		memory[16'h4380] <= 8'h70;
		memory[16'h4381] <= 8'h95;
		memory[16'h4382] <= 8'h82;
		memory[16'h4383] <= 8'h68;
		memory[16'h4384] <= 8'h87;
		memory[16'h4385] <= 8'hca;
		memory[16'h4386] <= 8'hfe;
		memory[16'h4387] <= 8'hcd;
		memory[16'h4388] <= 8'h9f;
		memory[16'h4389] <= 8'hda;
		memory[16'h438a] <= 8'h9;
		memory[16'h438b] <= 8'hdf;
		memory[16'h438c] <= 8'heb;
		memory[16'h438d] <= 8'h87;
		memory[16'h438e] <= 8'hc5;
		memory[16'h438f] <= 8'had;
		memory[16'h4390] <= 8'h6f;
		memory[16'h4391] <= 8'h45;
		memory[16'h4392] <= 8'h10;
		memory[16'h4393] <= 8'h86;
		memory[16'h4394] <= 8'h8;
		memory[16'h4395] <= 8'h4b;
		memory[16'h4396] <= 8'hef;
		memory[16'h4397] <= 8'h71;
		memory[16'h4398] <= 8'h54;
		memory[16'h4399] <= 8'h7;
		memory[16'h439a] <= 8'h7d;
		memory[16'h439b] <= 8'h3f;
		memory[16'h439c] <= 8'h12;
		memory[16'h439d] <= 8'h41;
		memory[16'h439e] <= 8'ha1;
		memory[16'h439f] <= 8'h82;
		memory[16'h43a0] <= 8'hd7;
		memory[16'h43a1] <= 8'h24;
		memory[16'h43a2] <= 8'hea;
		memory[16'h43a3] <= 8'h5e;
		memory[16'h43a4] <= 8'hee;
		memory[16'h43a5] <= 8'he8;
		memory[16'h43a6] <= 8'h2c;
		memory[16'h43a7] <= 8'h8e;
		memory[16'h43a8] <= 8'hc2;
		memory[16'h43a9] <= 8'h35;
		memory[16'h43aa] <= 8'h6d;
		memory[16'h43ab] <= 8'had;
		memory[16'h43ac] <= 8'hbd;
		memory[16'h43ad] <= 8'h33;
		memory[16'h43ae] <= 8'h5b;
		memory[16'h43af] <= 8'h2c;
		memory[16'h43b0] <= 8'h78;
		memory[16'h43b1] <= 8'h6b;
		memory[16'h43b2] <= 8'hb2;
		memory[16'h43b3] <= 8'h81;
		memory[16'h43b4] <= 8'hb6;
		memory[16'h43b5] <= 8'ha1;
		memory[16'h43b6] <= 8'hf2;
		memory[16'h43b7] <= 8'ha;
		memory[16'h43b8] <= 8'ha8;
		memory[16'h43b9] <= 8'h6f;
		memory[16'h43ba] <= 8'h49;
		memory[16'h43bb] <= 8'hba;
		memory[16'h43bc] <= 8'hb0;
		memory[16'h43bd] <= 8'heb;
		memory[16'h43be] <= 8'h3c;
		memory[16'h43bf] <= 8'h87;
		memory[16'h43c0] <= 8'hf;
		memory[16'h43c1] <= 8'h27;
		memory[16'h43c2] <= 8'he6;
		memory[16'h43c3] <= 8'hfd;
		memory[16'h43c4] <= 8'hf;
		memory[16'h43c5] <= 8'h12;
		memory[16'h43c6] <= 8'h8b;
		memory[16'h43c7] <= 8'hd2;
		memory[16'h43c8] <= 8'h47;
		memory[16'h43c9] <= 8'hf9;
		memory[16'h43ca] <= 8'h7f;
		memory[16'h43cb] <= 8'h4;
		memory[16'h43cc] <= 8'h2c;
		memory[16'h43cd] <= 8'hda;
		memory[16'h43ce] <= 8'h30;
		memory[16'h43cf] <= 8'ha4;
		memory[16'h43d0] <= 8'h45;
		memory[16'h43d1] <= 8'he2;
		memory[16'h43d2] <= 8'h25;
		memory[16'h43d3] <= 8'hfc;
		memory[16'h43d4] <= 8'h84;
		memory[16'h43d5] <= 8'h17;
		memory[16'h43d6] <= 8'h6;
		memory[16'h43d7] <= 8'h2c;
		memory[16'h43d8] <= 8'h86;
		memory[16'h43d9] <= 8'h50;
		memory[16'h43da] <= 8'he7;
		memory[16'h43db] <= 8'h37;
		memory[16'h43dc] <= 8'h3b;
		memory[16'h43dd] <= 8'h23;
		memory[16'h43de] <= 8'hbe;
		memory[16'h43df] <= 8'h4a;
		memory[16'h43e0] <= 8'h4a;
		memory[16'h43e1] <= 8'ha4;
		memory[16'h43e2] <= 8'h47;
		memory[16'h43e3] <= 8'h5a;
		memory[16'h43e4] <= 8'hb6;
		memory[16'h43e5] <= 8'hd3;
		memory[16'h43e6] <= 8'h2c;
		memory[16'h43e7] <= 8'hfe;
		memory[16'h43e8] <= 8'hcc;
		memory[16'h43e9] <= 8'hab;
		memory[16'h43ea] <= 8'h2;
		memory[16'h43eb] <= 8'hf8;
		memory[16'h43ec] <= 8'h86;
		memory[16'h43ed] <= 8'h33;
		memory[16'h43ee] <= 8'h9c;
		memory[16'h43ef] <= 8'hcb;
		memory[16'h43f0] <= 8'h15;
		memory[16'h43f1] <= 8'hc2;
		memory[16'h43f2] <= 8'hc7;
		memory[16'h43f3] <= 8'h99;
		memory[16'h43f4] <= 8'hd9;
		memory[16'h43f5] <= 8'hce;
		memory[16'h43f6] <= 8'hc6;
		memory[16'h43f7] <= 8'h60;
		memory[16'h43f8] <= 8'h1e;
		memory[16'h43f9] <= 8'had;
		memory[16'h43fa] <= 8'h97;
		memory[16'h43fb] <= 8'h59;
		memory[16'h43fc] <= 8'hd0;
		memory[16'h43fd] <= 8'h55;
		memory[16'h43fe] <= 8'ha3;
		memory[16'h43ff] <= 8'h1b;
		memory[16'h4400] <= 8'hfa;
		memory[16'h4401] <= 8'hea;
		memory[16'h4402] <= 8'h75;
		memory[16'h4403] <= 8'hb0;
		memory[16'h4404] <= 8'hbd;
		memory[16'h4405] <= 8'ha1;
		memory[16'h4406] <= 8'hae;
		memory[16'h4407] <= 8'h89;
		memory[16'h4408] <= 8'h4c;
		memory[16'h4409] <= 8'hb1;
		memory[16'h440a] <= 8'h81;
		memory[16'h440b] <= 8'hd2;
		memory[16'h440c] <= 8'he4;
		memory[16'h440d] <= 8'h1e;
		memory[16'h440e] <= 8'h9e;
		memory[16'h440f] <= 8'hf9;
		memory[16'h4410] <= 8'he0;
		memory[16'h4411] <= 8'h65;
		memory[16'h4412] <= 8'h93;
		memory[16'h4413] <= 8'hb9;
		memory[16'h4414] <= 8'h33;
		memory[16'h4415] <= 8'h59;
		memory[16'h4416] <= 8'h19;
		memory[16'h4417] <= 8'h51;
		memory[16'h4418] <= 8'h6;
		memory[16'h4419] <= 8'hb0;
		memory[16'h441a] <= 8'haa;
		memory[16'h441b] <= 8'hd6;
		memory[16'h441c] <= 8'h6;
		memory[16'h441d] <= 8'h4d;
		memory[16'h441e] <= 8'hf1;
		memory[16'h441f] <= 8'h0;
		memory[16'h4420] <= 8'h38;
		memory[16'h4421] <= 8'h66;
		memory[16'h4422] <= 8'hb0;
		memory[16'h4423] <= 8'hf5;
		memory[16'h4424] <= 8'h7;
		memory[16'h4425] <= 8'h5f;
		memory[16'h4426] <= 8'h7f;
		memory[16'h4427] <= 8'h54;
		memory[16'h4428] <= 8'h10;
		memory[16'h4429] <= 8'h0;
		memory[16'h442a] <= 8'h26;
		memory[16'h442b] <= 8'hf4;
		memory[16'h442c] <= 8'h1e;
		memory[16'h442d] <= 8'hc4;
		memory[16'h442e] <= 8'hed;
		memory[16'h442f] <= 8'hfe;
		memory[16'h4430] <= 8'h2a;
		memory[16'h4431] <= 8'h80;
		memory[16'h4432] <= 8'hb8;
		memory[16'h4433] <= 8'h5d;
		memory[16'h4434] <= 8'hd9;
		memory[16'h4435] <= 8'hd1;
		memory[16'h4436] <= 8'haf;
		memory[16'h4437] <= 8'hdf;
		memory[16'h4438] <= 8'h82;
		memory[16'h4439] <= 8'h59;
		memory[16'h443a] <= 8'hb6;
		memory[16'h443b] <= 8'h88;
		memory[16'h443c] <= 8'ha7;
		memory[16'h443d] <= 8'ha7;
		memory[16'h443e] <= 8'h88;
		memory[16'h443f] <= 8'hdf;
		memory[16'h4440] <= 8'he;
		memory[16'h4441] <= 8'h38;
		memory[16'h4442] <= 8'hd4;
		memory[16'h4443] <= 8'h15;
		memory[16'h4444] <= 8'h97;
		memory[16'h4445] <= 8'h53;
		memory[16'h4446] <= 8'h69;
		memory[16'h4447] <= 8'ha7;
		memory[16'h4448] <= 8'h54;
		memory[16'h4449] <= 8'h90;
		memory[16'h444a] <= 8'h9b;
		memory[16'h444b] <= 8'h72;
		memory[16'h444c] <= 8'h54;
		memory[16'h444d] <= 8'h89;
		memory[16'h444e] <= 8'h71;
		memory[16'h444f] <= 8'h7e;
		memory[16'h4450] <= 8'h9;
		memory[16'h4451] <= 8'h29;
		memory[16'h4452] <= 8'hdc;
		memory[16'h4453] <= 8'he3;
		memory[16'h4454] <= 8'hfa;
		memory[16'h4455] <= 8'h8b;
		memory[16'h4456] <= 8'hc2;
		memory[16'h4457] <= 8'h7c;
		memory[16'h4458] <= 8'he4;
		memory[16'h4459] <= 8'h78;
		memory[16'h445a] <= 8'h4;
		memory[16'h445b] <= 8'h8b;
		memory[16'h445c] <= 8'h20;
		memory[16'h445d] <= 8'h8c;
		memory[16'h445e] <= 8'h6a;
		memory[16'h445f] <= 8'h2e;
		memory[16'h4460] <= 8'hc5;
		memory[16'h4461] <= 8'h3f;
		memory[16'h4462] <= 8'h43;
		memory[16'h4463] <= 8'h5c;
		memory[16'h4464] <= 8'h92;
		memory[16'h4465] <= 8'had;
		memory[16'h4466] <= 8'h4;
		memory[16'h4467] <= 8'he6;
		memory[16'h4468] <= 8'h3d;
		memory[16'h4469] <= 8'h9f;
		memory[16'h446a] <= 8'h59;
		memory[16'h446b] <= 8'h91;
		memory[16'h446c] <= 8'h28;
		memory[16'h446d] <= 8'hca;
		memory[16'h446e] <= 8'h10;
		memory[16'h446f] <= 8'h32;
		memory[16'h4470] <= 8'hf3;
		memory[16'h4471] <= 8'hec;
		memory[16'h4472] <= 8'h15;
		memory[16'h4473] <= 8'hed;
		memory[16'h4474] <= 8'h77;
		memory[16'h4475] <= 8'hd7;
		memory[16'h4476] <= 8'h6a;
		memory[16'h4477] <= 8'h5b;
		memory[16'h4478] <= 8'h50;
		memory[16'h4479] <= 8'h6e;
		memory[16'h447a] <= 8'he7;
		memory[16'h447b] <= 8'h70;
		memory[16'h447c] <= 8'hfb;
		memory[16'h447d] <= 8'h51;
		memory[16'h447e] <= 8'h9e;
		memory[16'h447f] <= 8'hc0;
		memory[16'h4480] <= 8'h90;
		memory[16'h4481] <= 8'he1;
		memory[16'h4482] <= 8'h1c;
		memory[16'h4483] <= 8'h23;
		memory[16'h4484] <= 8'h8e;
		memory[16'h4485] <= 8'h20;
		memory[16'h4486] <= 8'h9;
		memory[16'h4487] <= 8'hcb;
		memory[16'h4488] <= 8'hc0;
		memory[16'h4489] <= 8'h62;
		memory[16'h448a] <= 8'h5d;
		memory[16'h448b] <= 8'he8;
		memory[16'h448c] <= 8'h2c;
		memory[16'h448d] <= 8'h6d;
		memory[16'h448e] <= 8'h1a;
		memory[16'h448f] <= 8'h1f;
		memory[16'h4490] <= 8'h59;
		memory[16'h4491] <= 8'h2f;
		memory[16'h4492] <= 8'hd;
		memory[16'h4493] <= 8'hd0;
		memory[16'h4494] <= 8'h7;
		memory[16'h4495] <= 8'h77;
		memory[16'h4496] <= 8'h2b;
		memory[16'h4497] <= 8'h57;
		memory[16'h4498] <= 8'he5;
		memory[16'h4499] <= 8'h12;
		memory[16'h449a] <= 8'hc7;
		memory[16'h449b] <= 8'he0;
		memory[16'h449c] <= 8'h64;
		memory[16'h449d] <= 8'h65;
		memory[16'h449e] <= 8'ha0;
		memory[16'h449f] <= 8'hf4;
		memory[16'h44a0] <= 8'h46;
		memory[16'h44a1] <= 8'hbd;
		memory[16'h44a2] <= 8'h17;
		memory[16'h44a3] <= 8'hd5;
		memory[16'h44a4] <= 8'hdd;
		memory[16'h44a5] <= 8'h21;
		memory[16'h44a6] <= 8'ha0;
		memory[16'h44a7] <= 8'h9d;
		memory[16'h44a8] <= 8'h83;
		memory[16'h44a9] <= 8'hfd;
		memory[16'h44aa] <= 8'h86;
		memory[16'h44ab] <= 8'hb0;
		memory[16'h44ac] <= 8'h6a;
		memory[16'h44ad] <= 8'ha0;
		memory[16'h44ae] <= 8'hcf;
		memory[16'h44af] <= 8'hc3;
		memory[16'h44b0] <= 8'hd0;
		memory[16'h44b1] <= 8'hdc;
		memory[16'h44b2] <= 8'h93;
		memory[16'h44b3] <= 8'hd7;
		memory[16'h44b4] <= 8'h53;
		memory[16'h44b5] <= 8'hbf;
		memory[16'h44b6] <= 8'h2e;
		memory[16'h44b7] <= 8'h39;
		memory[16'h44b8] <= 8'hd1;
		memory[16'h44b9] <= 8'hf5;
		memory[16'h44ba] <= 8'h19;
		memory[16'h44bb] <= 8'h35;
		memory[16'h44bc] <= 8'h5a;
		memory[16'h44bd] <= 8'hba;
		memory[16'h44be] <= 8'h2a;
		memory[16'h44bf] <= 8'ha0;
		memory[16'h44c0] <= 8'h77;
		memory[16'h44c1] <= 8'h41;
		memory[16'h44c2] <= 8'h75;
		memory[16'h44c3] <= 8'h54;
		memory[16'h44c4] <= 8'h62;
		memory[16'h44c5] <= 8'h16;
		memory[16'h44c6] <= 8'hf2;
		memory[16'h44c7] <= 8'he6;
		memory[16'h44c8] <= 8'h13;
		memory[16'h44c9] <= 8'h78;
		memory[16'h44ca] <= 8'h96;
		memory[16'h44cb] <= 8'h7e;
		memory[16'h44cc] <= 8'h18;
		memory[16'h44cd] <= 8'h65;
		memory[16'h44ce] <= 8'h41;
		memory[16'h44cf] <= 8'he8;
		memory[16'h44d0] <= 8'h42;
		memory[16'h44d1] <= 8'hd5;
		memory[16'h44d2] <= 8'hbf;
		memory[16'h44d3] <= 8'h95;
		memory[16'h44d4] <= 8'h94;
		memory[16'h44d5] <= 8'hed;
		memory[16'h44d6] <= 8'hce;
		memory[16'h44d7] <= 8'h65;
		memory[16'h44d8] <= 8'he2;
		memory[16'h44d9] <= 8'he8;
		memory[16'h44da] <= 8'h9b;
		memory[16'h44db] <= 8'h3c;
		memory[16'h44dc] <= 8'ha2;
		memory[16'h44dd] <= 8'hc5;
		memory[16'h44de] <= 8'hdd;
		memory[16'h44df] <= 8'h19;
		memory[16'h44e0] <= 8'h6;
		memory[16'h44e1] <= 8'h52;
		memory[16'h44e2] <= 8'h6d;
		memory[16'h44e3] <= 8'h69;
		memory[16'h44e4] <= 8'h68;
		memory[16'h44e5] <= 8'h5f;
		memory[16'h44e6] <= 8'h4f;
		memory[16'h44e7] <= 8'h7c;
		memory[16'h44e8] <= 8'hd7;
		memory[16'h44e9] <= 8'he5;
		memory[16'h44ea] <= 8'hfa;
		memory[16'h44eb] <= 8'hf0;
		memory[16'h44ec] <= 8'h4a;
		memory[16'h44ed] <= 8'h3b;
		memory[16'h44ee] <= 8'hd8;
		memory[16'h44ef] <= 8'h8c;
		memory[16'h44f0] <= 8'h10;
		memory[16'h44f1] <= 8'h98;
		memory[16'h44f2] <= 8'h22;
		memory[16'h44f3] <= 8'ha4;
		memory[16'h44f4] <= 8'h85;
		memory[16'h44f5] <= 8'hf0;
		memory[16'h44f6] <= 8'ha;
		memory[16'h44f7] <= 8'h68;
		memory[16'h44f8] <= 8'hd8;
		memory[16'h44f9] <= 8'ha5;
		memory[16'h44fa] <= 8'ha4;
		memory[16'h44fb] <= 8'h7a;
		memory[16'h44fc] <= 8'h6a;
		memory[16'h44fd] <= 8'h81;
		memory[16'h44fe] <= 8'h93;
		memory[16'h44ff] <= 8'h70;
		memory[16'h4500] <= 8'hd4;
		memory[16'h4501] <= 8'h1;
		memory[16'h4502] <= 8'hd9;
		memory[16'h4503] <= 8'h3c;
		memory[16'h4504] <= 8'h60;
		memory[16'h4505] <= 8'h28;
		memory[16'h4506] <= 8'hb8;
		memory[16'h4507] <= 8'h38;
		memory[16'h4508] <= 8'hd;
		memory[16'h4509] <= 8'hb2;
		memory[16'h450a] <= 8'h28;
		memory[16'h450b] <= 8'h58;
		memory[16'h450c] <= 8'hee;
		memory[16'h450d] <= 8'h0;
		memory[16'h450e] <= 8'he4;
		memory[16'h450f] <= 8'hfe;
		memory[16'h4510] <= 8'h98;
		memory[16'h4511] <= 8'h6;
		memory[16'h4512] <= 8'ha3;
		memory[16'h4513] <= 8'h1e;
		memory[16'h4514] <= 8'hf7;
		memory[16'h4515] <= 8'had;
		memory[16'h4516] <= 8'h86;
		memory[16'h4517] <= 8'hcf;
		memory[16'h4518] <= 8'h52;
		memory[16'h4519] <= 8'h2a;
		memory[16'h451a] <= 8'h4a;
		memory[16'h451b] <= 8'hbc;
		memory[16'h451c] <= 8'hac;
		memory[16'h451d] <= 8'hdd;
		memory[16'h451e] <= 8'h2c;
		memory[16'h451f] <= 8'h80;
		memory[16'h4520] <= 8'hde;
		memory[16'h4521] <= 8'h6;
		memory[16'h4522] <= 8'hbc;
		memory[16'h4523] <= 8'h3f;
		memory[16'h4524] <= 8'h2e;
		memory[16'h4525] <= 8'h75;
		memory[16'h4526] <= 8'h77;
		memory[16'h4527] <= 8'h3c;
		memory[16'h4528] <= 8'h27;
		memory[16'h4529] <= 8'h9f;
		memory[16'h452a] <= 8'h94;
		memory[16'h452b] <= 8'h15;
		memory[16'h452c] <= 8'h9f;
		memory[16'h452d] <= 8'h78;
		memory[16'h452e] <= 8'h14;
		memory[16'h452f] <= 8'h38;
		memory[16'h4530] <= 8'h7f;
		memory[16'h4531] <= 8'hb7;
		memory[16'h4532] <= 8'h56;
		memory[16'h4533] <= 8'h76;
		memory[16'h4534] <= 8'h64;
		memory[16'h4535] <= 8'hdc;
		memory[16'h4536] <= 8'h45;
		memory[16'h4537] <= 8'hb6;
		memory[16'h4538] <= 8'h6;
		memory[16'h4539] <= 8'h8f;
		memory[16'h453a] <= 8'h72;
		memory[16'h453b] <= 8'hb2;
		memory[16'h453c] <= 8'h6d;
		memory[16'h453d] <= 8'h9e;
		memory[16'h453e] <= 8'h32;
		memory[16'h453f] <= 8'h4b;
		memory[16'h4540] <= 8'ha4;
		memory[16'h4541] <= 8'hef;
		memory[16'h4542] <= 8'h8a;
		memory[16'h4543] <= 8'hd3;
		memory[16'h4544] <= 8'h64;
		memory[16'h4545] <= 8'h1;
		memory[16'h4546] <= 8'hf;
		memory[16'h4547] <= 8'h8b;
		memory[16'h4548] <= 8'ha0;
		memory[16'h4549] <= 8'ha3;
		memory[16'h454a] <= 8'ha1;
		memory[16'h454b] <= 8'h40;
		memory[16'h454c] <= 8'h1b;
		memory[16'h454d] <= 8'hb5;
		memory[16'h454e] <= 8'h78;
		memory[16'h454f] <= 8'h9a;
		memory[16'h4550] <= 8'h6c;
		memory[16'h4551] <= 8'hce;
		memory[16'h4552] <= 8'h10;
		memory[16'h4553] <= 8'hd0;
		memory[16'h4554] <= 8'haa;
		memory[16'h4555] <= 8'h56;
		memory[16'h4556] <= 8'h86;
		memory[16'h4557] <= 8'hb0;
		memory[16'h4558] <= 8'he5;
		memory[16'h4559] <= 8'hf8;
		memory[16'h455a] <= 8'h63;
		memory[16'h455b] <= 8'h52;
		memory[16'h455c] <= 8'h96;
		memory[16'h455d] <= 8'h95;
		memory[16'h455e] <= 8'h9e;
		memory[16'h455f] <= 8'h3b;
		memory[16'h4560] <= 8'h84;
		memory[16'h4561] <= 8'h28;
		memory[16'h4562] <= 8'he;
		memory[16'h4563] <= 8'he8;
		memory[16'h4564] <= 8'h2a;
		memory[16'h4565] <= 8'h1d;
		memory[16'h4566] <= 8'h74;
		memory[16'h4567] <= 8'hca;
		memory[16'h4568] <= 8'hc0;
		memory[16'h4569] <= 8'h15;
		memory[16'h456a] <= 8'ha;
		memory[16'h456b] <= 8'hdb;
		memory[16'h456c] <= 8'hca;
		memory[16'h456d] <= 8'h82;
		memory[16'h456e] <= 8'h76;
		memory[16'h456f] <= 8'h36;
		memory[16'h4570] <= 8'h50;
		memory[16'h4571] <= 8'h86;
		memory[16'h4572] <= 8'h6;
		memory[16'h4573] <= 8'hfa;
		memory[16'h4574] <= 8'hdc;
		memory[16'h4575] <= 8'h8c;
		memory[16'h4576] <= 8'hab;
		memory[16'h4577] <= 8'hc2;
		memory[16'h4578] <= 8'h84;
		memory[16'h4579] <= 8'he;
		memory[16'h457a] <= 8'h14;
		memory[16'h457b] <= 8'h1a;
		memory[16'h457c] <= 8'ha3;
		memory[16'h457d] <= 8'hb2;
		memory[16'h457e] <= 8'h55;
		memory[16'h457f] <= 8'h28;
		memory[16'h4580] <= 8'hdb;
		memory[16'h4581] <= 8'h63;
		memory[16'h4582] <= 8'h10;
		memory[16'h4583] <= 8'h5;
		memory[16'h4584] <= 8'h80;
		memory[16'h4585] <= 8'h84;
		memory[16'h4586] <= 8'hcf;
		memory[16'h4587] <= 8'h40;
		memory[16'h4588] <= 8'h99;
		memory[16'h4589] <= 8'hda;
		memory[16'h458a] <= 8'h1c;
		memory[16'h458b] <= 8'h63;
		memory[16'h458c] <= 8'h5c;
		memory[16'h458d] <= 8'h92;
		memory[16'h458e] <= 8'h99;
		memory[16'h458f] <= 8'had;
		memory[16'h4590] <= 8'h18;
		memory[16'h4591] <= 8'h9f;
		memory[16'h4592] <= 8'ha7;
		memory[16'h4593] <= 8'hf5;
		memory[16'h4594] <= 8'h2b;
		memory[16'h4595] <= 8'h52;
		memory[16'h4596] <= 8'hb7;
		memory[16'h4597] <= 8'haf;
		memory[16'h4598] <= 8'h60;
		memory[16'h4599] <= 8'hcb;
		memory[16'h459a] <= 8'hca;
		memory[16'h459b] <= 8'h4;
		memory[16'h459c] <= 8'h7e;
		memory[16'h459d] <= 8'h1f;
		memory[16'h459e] <= 8'h2c;
		memory[16'h459f] <= 8'h59;
		memory[16'h45a0] <= 8'h83;
		memory[16'h45a1] <= 8'h3c;
		memory[16'h45a2] <= 8'h5e;
		memory[16'h45a3] <= 8'h3;
		memory[16'h45a4] <= 8'hc1;
		memory[16'h45a5] <= 8'h2d;
		memory[16'h45a6] <= 8'h44;
		memory[16'h45a7] <= 8'h5a;
		memory[16'h45a8] <= 8'h7;
		memory[16'h45a9] <= 8'h60;
		memory[16'h45aa] <= 8'hbe;
		memory[16'h45ab] <= 8'h64;
		memory[16'h45ac] <= 8'hf2;
		memory[16'h45ad] <= 8'h57;
		memory[16'h45ae] <= 8'h11;
		memory[16'h45af] <= 8'ha;
		memory[16'h45b0] <= 8'hf7;
		memory[16'h45b1] <= 8'hb8;
		memory[16'h45b2] <= 8'hff;
		memory[16'h45b3] <= 8'h22;
		memory[16'h45b4] <= 8'hb;
		memory[16'h45b5] <= 8'hb6;
		memory[16'h45b6] <= 8'hd2;
		memory[16'h45b7] <= 8'h6b;
		memory[16'h45b8] <= 8'h82;
		memory[16'h45b9] <= 8'h9c;
		memory[16'h45ba] <= 8'h6f;
		memory[16'h45bb] <= 8'h0;
		memory[16'h45bc] <= 8'hbb;
		memory[16'h45bd] <= 8'h9b;
		memory[16'h45be] <= 8'h59;
		memory[16'h45bf] <= 8'h3e;
		memory[16'h45c0] <= 8'hd8;
		memory[16'h45c1] <= 8'hb7;
		memory[16'h45c2] <= 8'h42;
		memory[16'h45c3] <= 8'h99;
		memory[16'h45c4] <= 8'he4;
		memory[16'h45c5] <= 8'h86;
		memory[16'h45c6] <= 8'hf3;
		memory[16'h45c7] <= 8'hec;
		memory[16'h45c8] <= 8'he6;
		memory[16'h45c9] <= 8'hb1;
		memory[16'h45ca] <= 8'h50;
		memory[16'h45cb] <= 8'hd8;
		memory[16'h45cc] <= 8'h9;
		memory[16'h45cd] <= 8'h61;
		memory[16'h45ce] <= 8'he2;
		memory[16'h45cf] <= 8'h0;
		memory[16'h45d0] <= 8'h19;
		memory[16'h45d1] <= 8'he2;
		memory[16'h45d2] <= 8'h22;
		memory[16'h45d3] <= 8'h24;
		memory[16'h45d4] <= 8'h98;
		memory[16'h45d5] <= 8'hf4;
		memory[16'h45d6] <= 8'h90;
		memory[16'h45d7] <= 8'h1a;
		memory[16'h45d8] <= 8'h90;
		memory[16'h45d9] <= 8'hff;
		memory[16'h45da] <= 8'h1a;
		memory[16'h45db] <= 8'h4c;
		memory[16'h45dc] <= 8'h9b;
		memory[16'h45dd] <= 8'h73;
		memory[16'h45de] <= 8'h8a;
		memory[16'h45df] <= 8'h73;
		memory[16'h45e0] <= 8'h2a;
		memory[16'h45e1] <= 8'hcc;
		memory[16'h45e2] <= 8'hc;
		memory[16'h45e3] <= 8'hf;
		memory[16'h45e4] <= 8'h52;
		memory[16'h45e5] <= 8'hff;
		memory[16'h45e6] <= 8'hfb;
		memory[16'h45e7] <= 8'h38;
		memory[16'h45e8] <= 8'hb1;
		memory[16'h45e9] <= 8'h4b;
		memory[16'h45ea] <= 8'h10;
		memory[16'h45eb] <= 8'hba;
		memory[16'h45ec] <= 8'hac;
		memory[16'h45ed] <= 8'hf3;
		memory[16'h45ee] <= 8'hba;
		memory[16'h45ef] <= 8'hc5;
		memory[16'h45f0] <= 8'hd5;
		memory[16'h45f1] <= 8'hdc;
		memory[16'h45f2] <= 8'hea;
		memory[16'h45f3] <= 8'h6d;
		memory[16'h45f4] <= 8'hd1;
		memory[16'h45f5] <= 8'h7a;
		memory[16'h45f6] <= 8'h88;
		memory[16'h45f7] <= 8'h61;
		memory[16'h45f8] <= 8'h79;
		memory[16'h45f9] <= 8'ha2;
		memory[16'h45fa] <= 8'had;
		memory[16'h45fb] <= 8'h14;
		memory[16'h45fc] <= 8'h16;
		memory[16'h45fd] <= 8'h38;
		memory[16'h45fe] <= 8'h87;
		memory[16'h45ff] <= 8'h40;
		memory[16'h4600] <= 8'h4;
		memory[16'h4601] <= 8'h93;
		memory[16'h4602] <= 8'h4f;
		memory[16'h4603] <= 8'h57;
		memory[16'h4604] <= 8'h93;
		memory[16'h4605] <= 8'h4a;
		memory[16'h4606] <= 8'h8f;
		memory[16'h4607] <= 8'h44;
		memory[16'h4608] <= 8'h95;
		memory[16'h4609] <= 8'ha0;
		memory[16'h460a] <= 8'hfe;
		memory[16'h460b] <= 8'h41;
		memory[16'h460c] <= 8'h93;
		memory[16'h460d] <= 8'hb8;
		memory[16'h460e] <= 8'h7;
		memory[16'h460f] <= 8'h68;
		memory[16'h4610] <= 8'h94;
		memory[16'h4611] <= 8'hf1;
		memory[16'h4612] <= 8'hd5;
		memory[16'h4613] <= 8'h65;
		memory[16'h4614] <= 8'h6b;
		memory[16'h4615] <= 8'h5d;
		memory[16'h4616] <= 8'hc7;
		memory[16'h4617] <= 8'he4;
		memory[16'h4618] <= 8'h0;
		memory[16'h4619] <= 8'h74;
		memory[16'h461a] <= 8'hf9;
		memory[16'h461b] <= 8'h16;
		memory[16'h461c] <= 8'hac;
		memory[16'h461d] <= 8'h80;
		memory[16'h461e] <= 8'h56;
		memory[16'h461f] <= 8'hb1;
		memory[16'h4620] <= 8'h14;
		memory[16'h4621] <= 8'ha6;
		memory[16'h4622] <= 8'h8;
		memory[16'h4623] <= 8'ha7;
		memory[16'h4624] <= 8'hf0;
		memory[16'h4625] <= 8'h97;
		memory[16'h4626] <= 8'heb;
		memory[16'h4627] <= 8'h86;
		memory[16'h4628] <= 8'h37;
		memory[16'h4629] <= 8'he9;
		memory[16'h462a] <= 8'hc7;
		memory[16'h462b] <= 8'hca;
		memory[16'h462c] <= 8'ha1;
		memory[16'h462d] <= 8'hce;
		memory[16'h462e] <= 8'h32;
		memory[16'h462f] <= 8'h35;
		memory[16'h4630] <= 8'hbf;
		memory[16'h4631] <= 8'h8;
		memory[16'h4632] <= 8'h9b;
		memory[16'h4633] <= 8'h2a;
		memory[16'h4634] <= 8'h65;
		memory[16'h4635] <= 8'h62;
		memory[16'h4636] <= 8'hf;
		memory[16'h4637] <= 8'h65;
		memory[16'h4638] <= 8'hd6;
		memory[16'h4639] <= 8'h8;
		memory[16'h463a] <= 8'h7b;
		memory[16'h463b] <= 8'h83;
		memory[16'h463c] <= 8'h88;
		memory[16'h463d] <= 8'hd2;
		memory[16'h463e] <= 8'h34;
		memory[16'h463f] <= 8'h9c;
		memory[16'h4640] <= 8'h78;
		memory[16'h4641] <= 8'h3c;
		memory[16'h4642] <= 8'h43;
		memory[16'h4643] <= 8'h68;
		memory[16'h4644] <= 8'hd3;
		memory[16'h4645] <= 8'h2e;
		memory[16'h4646] <= 8'hee;
		memory[16'h4647] <= 8'hb;
		memory[16'h4648] <= 8'h17;
		memory[16'h4649] <= 8'hb6;
		memory[16'h464a] <= 8'hd5;
		memory[16'h464b] <= 8'hb8;
		memory[16'h464c] <= 8'h84;
		memory[16'h464d] <= 8'h8;
		memory[16'h464e] <= 8'hee;
		memory[16'h464f] <= 8'h44;
		memory[16'h4650] <= 8'h10;
		memory[16'h4651] <= 8'h89;
		memory[16'h4652] <= 8'h6e;
		memory[16'h4653] <= 8'h75;
		memory[16'h4654] <= 8'heb;
		memory[16'h4655] <= 8'h7d;
		memory[16'h4656] <= 8'hdb;
		memory[16'h4657] <= 8'hc1;
		memory[16'h4658] <= 8'h85;
		memory[16'h4659] <= 8'h56;
		memory[16'h465a] <= 8'h44;
		memory[16'h465b] <= 8'he;
		memory[16'h465c] <= 8'h28;
		memory[16'h465d] <= 8'h78;
		memory[16'h465e] <= 8'haa;
		memory[16'h465f] <= 8'ha0;
		memory[16'h4660] <= 8'hb4;
		memory[16'h4661] <= 8'hee;
		memory[16'h4662] <= 8'h9;
		memory[16'h4663] <= 8'h88;
		memory[16'h4664] <= 8'h1c;
		memory[16'h4665] <= 8'hf7;
		memory[16'h4666] <= 8'h93;
		memory[16'h4667] <= 8'h34;
		memory[16'h4668] <= 8'had;
		memory[16'h4669] <= 8'h68;
		memory[16'h466a] <= 8'hec;
		memory[16'h466b] <= 8'h32;
		memory[16'h466c] <= 8'h70;
		memory[16'h466d] <= 8'hda;
		memory[16'h466e] <= 8'h76;
		memory[16'h466f] <= 8'h80;
		memory[16'h4670] <= 8'h63;
		memory[16'h4671] <= 8'he4;
		memory[16'h4672] <= 8'hf6;
		memory[16'h4673] <= 8'h4e;
		memory[16'h4674] <= 8'h62;
		memory[16'h4675] <= 8'hd1;
		memory[16'h4676] <= 8'h10;
		memory[16'h4677] <= 8'he7;
		memory[16'h4678] <= 8'h27;
		memory[16'h4679] <= 8'h54;
		memory[16'h467a] <= 8'hf5;
		memory[16'h467b] <= 8'h50;
		memory[16'h467c] <= 8'hcd;
		memory[16'h467d] <= 8'ha0;
		memory[16'h467e] <= 8'hf0;
		memory[16'h467f] <= 8'h81;
		memory[16'h4680] <= 8'h8e;
		memory[16'h4681] <= 8'hf9;
		memory[16'h4682] <= 8'h9;
		memory[16'h4683] <= 8'haa;
		memory[16'h4684] <= 8'hf1;
		memory[16'h4685] <= 8'h9c;
		memory[16'h4686] <= 8'hde;
		memory[16'h4687] <= 8'h9e;
		memory[16'h4688] <= 8'h5;
		memory[16'h4689] <= 8'hcb;
		memory[16'h468a] <= 8'hd0;
		memory[16'h468b] <= 8'h75;
		memory[16'h468c] <= 8'ha5;
		memory[16'h468d] <= 8'h46;
		memory[16'h468e] <= 8'hf6;
		memory[16'h468f] <= 8'h9;
		memory[16'h4690] <= 8'h2b;
		memory[16'h4691] <= 8'hec;
		memory[16'h4692] <= 8'h57;
		memory[16'h4693] <= 8'h8d;
		memory[16'h4694] <= 8'hbd;
		memory[16'h4695] <= 8'h67;
		memory[16'h4696] <= 8'h74;
		memory[16'h4697] <= 8'he4;
		memory[16'h4698] <= 8'hbc;
		memory[16'h4699] <= 8'h6a;
		memory[16'h469a] <= 8'h34;
		memory[16'h469b] <= 8'h89;
		memory[16'h469c] <= 8'ha;
		memory[16'h469d] <= 8'h25;
		memory[16'h469e] <= 8'ha;
		memory[16'h469f] <= 8'h98;
		memory[16'h46a0] <= 8'h1e;
		memory[16'h46a1] <= 8'h14;
		memory[16'h46a2] <= 8'h42;
		memory[16'h46a3] <= 8'hf;
		memory[16'h46a4] <= 8'hb0;
		memory[16'h46a5] <= 8'h21;
		memory[16'h46a6] <= 8'hae;
		memory[16'h46a7] <= 8'hb5;
		memory[16'h46a8] <= 8'hec;
		memory[16'h46a9] <= 8'h7e;
		memory[16'h46aa] <= 8'h2b;
		memory[16'h46ab] <= 8'h91;
		memory[16'h46ac] <= 8'hc5;
		memory[16'h46ad] <= 8'h21;
		memory[16'h46ae] <= 8'h9a;
		memory[16'h46af] <= 8'hf0;
		memory[16'h46b0] <= 8'hd;
		memory[16'h46b1] <= 8'hf2;
		memory[16'h46b2] <= 8'h7d;
		memory[16'h46b3] <= 8'hca;
		memory[16'h46b4] <= 8'h59;
		memory[16'h46b5] <= 8'hf1;
		memory[16'h46b6] <= 8'hae;
		memory[16'h46b7] <= 8'h15;
		memory[16'h46b8] <= 8'h5b;
		memory[16'h46b9] <= 8'he3;
		memory[16'h46ba] <= 8'h9e;
		memory[16'h46bb] <= 8'h65;
		memory[16'h46bc] <= 8'h8;
		memory[16'h46bd] <= 8'ha9;
		memory[16'h46be] <= 8'hfd;
		memory[16'h46bf] <= 8'h26;
		memory[16'h46c0] <= 8'hbd;
		memory[16'h46c1] <= 8'h40;
		memory[16'h46c2] <= 8'h36;
		memory[16'h46c3] <= 8'h6d;
		memory[16'h46c4] <= 8'h61;
		memory[16'h46c5] <= 8'he4;
		memory[16'h46c6] <= 8'h23;
		memory[16'h46c7] <= 8'h4d;
		memory[16'h46c8] <= 8'h62;
		memory[16'h46c9] <= 8'h4e;
		memory[16'h46ca] <= 8'hde;
		memory[16'h46cb] <= 8'h27;
		memory[16'h46cc] <= 8'h6f;
		memory[16'h46cd] <= 8'h79;
		memory[16'h46ce] <= 8'h17;
		memory[16'h46cf] <= 8'h7c;
		memory[16'h46d0] <= 8'h6b;
		memory[16'h46d1] <= 8'h94;
		memory[16'h46d2] <= 8'h46;
		memory[16'h46d3] <= 8'hc4;
		memory[16'h46d4] <= 8'h86;
		memory[16'h46d5] <= 8'hf4;
		memory[16'h46d6] <= 8'hda;
		memory[16'h46d7] <= 8'he1;
		memory[16'h46d8] <= 8'hd7;
		memory[16'h46d9] <= 8'h78;
		memory[16'h46da] <= 8'h47;
		memory[16'h46db] <= 8'hdf;
		memory[16'h46dc] <= 8'h21;
		memory[16'h46dd] <= 8'h44;
		memory[16'h46de] <= 8'h6;
		memory[16'h46df] <= 8'hde;
		memory[16'h46e0] <= 8'h84;
		memory[16'h46e1] <= 8'h3c;
		memory[16'h46e2] <= 8'h4c;
		memory[16'h46e3] <= 8'he5;
		memory[16'h46e4] <= 8'h20;
		memory[16'h46e5] <= 8'h6f;
		memory[16'h46e6] <= 8'h32;
		memory[16'h46e7] <= 8'h82;
		memory[16'h46e8] <= 8'hbd;
		memory[16'h46e9] <= 8'h11;
		memory[16'h46ea] <= 8'haa;
		memory[16'h46eb] <= 8'h2c;
		memory[16'h46ec] <= 8'h8a;
		memory[16'h46ed] <= 8'hc1;
		memory[16'h46ee] <= 8'ha8;
		memory[16'h46ef] <= 8'hf5;
		memory[16'h46f0] <= 8'h56;
		memory[16'h46f1] <= 8'hee;
		memory[16'h46f2] <= 8'hb9;
		memory[16'h46f3] <= 8'hdc;
		memory[16'h46f4] <= 8'he2;
		memory[16'h46f5] <= 8'h93;
		memory[16'h46f6] <= 8'hbd;
		memory[16'h46f7] <= 8'hba;
		memory[16'h46f8] <= 8'hc;
		memory[16'h46f9] <= 8'h4;
		memory[16'h46fa] <= 8'h99;
		memory[16'h46fb] <= 8'h2d;
		memory[16'h46fc] <= 8'h49;
		memory[16'h46fd] <= 8'h9f;
		memory[16'h46fe] <= 8'hc;
		memory[16'h46ff] <= 8'hcd;
		memory[16'h4700] <= 8'hdb;
		memory[16'h4701] <= 8'h58;
		memory[16'h4702] <= 8'hb3;
		memory[16'h4703] <= 8'hfb;
		memory[16'h4704] <= 8'hc7;
		memory[16'h4705] <= 8'he5;
		memory[16'h4706] <= 8'h7e;
		memory[16'h4707] <= 8'h84;
		memory[16'h4708] <= 8'hf6;
		memory[16'h4709] <= 8'h28;
		memory[16'h470a] <= 8'hb0;
		memory[16'h470b] <= 8'h80;
		memory[16'h470c] <= 8'he9;
		memory[16'h470d] <= 8'h58;
		memory[16'h470e] <= 8'h75;
		memory[16'h470f] <= 8'h3f;
		memory[16'h4710] <= 8'h46;
		memory[16'h4711] <= 8'h2f;
		memory[16'h4712] <= 8'h1b;
		memory[16'h4713] <= 8'h28;
		memory[16'h4714] <= 8'hc2;
		memory[16'h4715] <= 8'hd9;
		memory[16'h4716] <= 8'he2;
		memory[16'h4717] <= 8'hce;
		memory[16'h4718] <= 8'hdd;
		memory[16'h4719] <= 8'h7c;
		memory[16'h471a] <= 8'hfc;
		memory[16'h471b] <= 8'h26;
		memory[16'h471c] <= 8'h1b;
		memory[16'h471d] <= 8'h8;
		memory[16'h471e] <= 8'hf4;
		memory[16'h471f] <= 8'hf7;
		memory[16'h4720] <= 8'h60;
		memory[16'h4721] <= 8'ha7;
		memory[16'h4722] <= 8'hf2;
		memory[16'h4723] <= 8'h27;
		memory[16'h4724] <= 8'h8c;
		memory[16'h4725] <= 8'h70;
		memory[16'h4726] <= 8'hab;
		memory[16'h4727] <= 8'h83;
		memory[16'h4728] <= 8'h98;
		memory[16'h4729] <= 8'h5b;
		memory[16'h472a] <= 8'h3;
		memory[16'h472b] <= 8'h82;
		memory[16'h472c] <= 8'hb3;
		memory[16'h472d] <= 8'h79;
		memory[16'h472e] <= 8'hc1;
		memory[16'h472f] <= 8'hf9;
		memory[16'h4730] <= 8'ha8;
		memory[16'h4731] <= 8'hdd;
		memory[16'h4732] <= 8'h21;
		memory[16'h4733] <= 8'h6a;
		memory[16'h4734] <= 8'hb6;
		memory[16'h4735] <= 8'h4;
		memory[16'h4736] <= 8'h39;
		memory[16'h4737] <= 8'h93;
		memory[16'h4738] <= 8'h80;
		memory[16'h4739] <= 8'h35;
		memory[16'h473a] <= 8'hba;
		memory[16'h473b] <= 8'h9b;
		memory[16'h473c] <= 8'h3d;
		memory[16'h473d] <= 8'hae;
		memory[16'h473e] <= 8'h92;
		memory[16'h473f] <= 8'h9d;
		memory[16'h4740] <= 8'h55;
		memory[16'h4741] <= 8'h85;
		memory[16'h4742] <= 8'hc4;
		memory[16'h4743] <= 8'he1;
		memory[16'h4744] <= 8'hf5;
		memory[16'h4745] <= 8'h6f;
		memory[16'h4746] <= 8'h64;
		memory[16'h4747] <= 8'h8e;
		memory[16'h4748] <= 8'hca;
		memory[16'h4749] <= 8'h68;
		memory[16'h474a] <= 8'h10;
		memory[16'h474b] <= 8'h7d;
		memory[16'h474c] <= 8'he1;
		memory[16'h474d] <= 8'hd1;
		memory[16'h474e] <= 8'h76;
		memory[16'h474f] <= 8'h89;
		memory[16'h4750] <= 8'hae;
		memory[16'h4751] <= 8'h97;
		memory[16'h4752] <= 8'hf3;
		memory[16'h4753] <= 8'h64;
		memory[16'h4754] <= 8'h9b;
		memory[16'h4755] <= 8'h2c;
		memory[16'h4756] <= 8'hf8;
		memory[16'h4757] <= 8'h1b;
		memory[16'h4758] <= 8'h61;
		memory[16'h4759] <= 8'hb2;
		memory[16'h475a] <= 8'hb7;
		memory[16'h475b] <= 8'h9e;
		memory[16'h475c] <= 8'h60;
		memory[16'h475d] <= 8'h49;
		memory[16'h475e] <= 8'h3b;
		memory[16'h475f] <= 8'hb5;
		memory[16'h4760] <= 8'hce;
		memory[16'h4761] <= 8'hff;
		memory[16'h4762] <= 8'h96;
		memory[16'h4763] <= 8'hc4;
		memory[16'h4764] <= 8'h6e;
		memory[16'h4765] <= 8'hfb;
		memory[16'h4766] <= 8'h52;
		memory[16'h4767] <= 8'h38;
		memory[16'h4768] <= 8'h63;
		memory[16'h4769] <= 8'h62;
		memory[16'h476a] <= 8'hb5;
		memory[16'h476b] <= 8'h44;
		memory[16'h476c] <= 8'h33;
		memory[16'h476d] <= 8'h2b;
		memory[16'h476e] <= 8'hcd;
		memory[16'h476f] <= 8'he2;
		memory[16'h4770] <= 8'hc3;
		memory[16'h4771] <= 8'hc0;
		memory[16'h4772] <= 8'h46;
		memory[16'h4773] <= 8'h5e;
		memory[16'h4774] <= 8'hed;
		memory[16'h4775] <= 8'h3e;
		memory[16'h4776] <= 8'h7a;
		memory[16'h4777] <= 8'h4e;
		memory[16'h4778] <= 8'hf0;
		memory[16'h4779] <= 8'h31;
		memory[16'h477a] <= 8'hed;
		memory[16'h477b] <= 8'h50;
		memory[16'h477c] <= 8'h7a;
		memory[16'h477d] <= 8'h28;
		memory[16'h477e] <= 8'h5;
		memory[16'h477f] <= 8'h49;
		memory[16'h4780] <= 8'h28;
		memory[16'h4781] <= 8'h9c;
		memory[16'h4782] <= 8'hd;
		memory[16'h4783] <= 8'h96;
		memory[16'h4784] <= 8'h97;
		memory[16'h4785] <= 8'h5f;
		memory[16'h4786] <= 8'hcf;
		memory[16'h4787] <= 8'hfa;
		memory[16'h4788] <= 8'hc1;
		memory[16'h4789] <= 8'h84;
		memory[16'h478a] <= 8'h3e;
		memory[16'h478b] <= 8'hf4;
		memory[16'h478c] <= 8'hb0;
		memory[16'h478d] <= 8'hb;
		memory[16'h478e] <= 8'hd6;
		memory[16'h478f] <= 8'h73;
		memory[16'h4790] <= 8'hcb;
		memory[16'h4791] <= 8'h1d;
		memory[16'h4792] <= 8'hd1;
		memory[16'h4793] <= 8'hb8;
		memory[16'h4794] <= 8'h5b;
		memory[16'h4795] <= 8'h4b;
		memory[16'h4796] <= 8'h7;
		memory[16'h4797] <= 8'h4c;
		memory[16'h4798] <= 8'h7c;
		memory[16'h4799] <= 8'hf4;
		memory[16'h479a] <= 8'h9c;
		memory[16'h479b] <= 8'hf7;
		memory[16'h479c] <= 8'h1c;
		memory[16'h479d] <= 8'ha2;
		memory[16'h479e] <= 8'h40;
		memory[16'h479f] <= 8'h44;
		memory[16'h47a0] <= 8'h3e;
		memory[16'h47a1] <= 8'h4d;
		memory[16'h47a2] <= 8'hdb;
		memory[16'h47a3] <= 8'hd5;
		memory[16'h47a4] <= 8'hac;
		memory[16'h47a5] <= 8'haa;
		memory[16'h47a6] <= 8'hcf;
		memory[16'h47a7] <= 8'h6d;
		memory[16'h47a8] <= 8'h2e;
		memory[16'h47a9] <= 8'hd;
		memory[16'h47aa] <= 8'h61;
		memory[16'h47ab] <= 8'hde;
		memory[16'h47ac] <= 8'h18;
		memory[16'h47ad] <= 8'h38;
		memory[16'h47ae] <= 8'h51;
		memory[16'h47af] <= 8'he3;
		memory[16'h47b0] <= 8'h55;
		memory[16'h47b1] <= 8'h23;
		memory[16'h47b2] <= 8'h9c;
		memory[16'h47b3] <= 8'hb0;
		memory[16'h47b4] <= 8'h6e;
		memory[16'h47b5] <= 8'ha3;
		memory[16'h47b6] <= 8'hfc;
		memory[16'h47b7] <= 8'heb;
		memory[16'h47b8] <= 8'h97;
		memory[16'h47b9] <= 8'h99;
		memory[16'h47ba] <= 8'he2;
		memory[16'h47bb] <= 8'hb3;
		memory[16'h47bc] <= 8'h3b;
		memory[16'h47bd] <= 8'h22;
		memory[16'h47be] <= 8'hf8;
		memory[16'h47bf] <= 8'h79;
		memory[16'h47c0] <= 8'h6f;
		memory[16'h47c1] <= 8'hd3;
		memory[16'h47c2] <= 8'h4e;
		memory[16'h47c3] <= 8'h1b;
		memory[16'h47c4] <= 8'h7d;
		memory[16'h47c5] <= 8'h1d;
		memory[16'h47c6] <= 8'h88;
		memory[16'h47c7] <= 8'hab;
		memory[16'h47c8] <= 8'h2a;
		memory[16'h47c9] <= 8'he9;
		memory[16'h47ca] <= 8'h8a;
		memory[16'h47cb] <= 8'h42;
		memory[16'h47cc] <= 8'h21;
		memory[16'h47cd] <= 8'hdb;
		memory[16'h47ce] <= 8'h25;
		memory[16'h47cf] <= 8'h76;
		memory[16'h47d0] <= 8'hfe;
		memory[16'h47d1] <= 8'hc1;
		memory[16'h47d2] <= 8'h27;
		memory[16'h47d3] <= 8'h6d;
		memory[16'h47d4] <= 8'h64;
		memory[16'h47d5] <= 8'h23;
		memory[16'h47d6] <= 8'h58;
		memory[16'h47d7] <= 8'hfb;
		memory[16'h47d8] <= 8'hbc;
		memory[16'h47d9] <= 8'h3a;
		memory[16'h47da] <= 8'haf;
		memory[16'h47db] <= 8'hf7;
		memory[16'h47dc] <= 8'h5c;
		memory[16'h47dd] <= 8'ha7;
		memory[16'h47de] <= 8'h70;
		memory[16'h47df] <= 8'hcb;
		memory[16'h47e0] <= 8'h7a;
		memory[16'h47e1] <= 8'hbe;
		memory[16'h47e2] <= 8'he6;
		memory[16'h47e3] <= 8'hf7;
		memory[16'h47e4] <= 8'hdb;
		memory[16'h47e5] <= 8'h6e;
		memory[16'h47e6] <= 8'ha2;
		memory[16'h47e7] <= 8'h5;
		memory[16'h47e8] <= 8'h57;
		memory[16'h47e9] <= 8'h2c;
		memory[16'h47ea] <= 8'h47;
		memory[16'h47eb] <= 8'h79;
		memory[16'h47ec] <= 8'h8;
		memory[16'h47ed] <= 8'h6d;
		memory[16'h47ee] <= 8'hef;
		memory[16'h47ef] <= 8'h6;
		memory[16'h47f0] <= 8'h2e;
		memory[16'h47f1] <= 8'h16;
		memory[16'h47f2] <= 8'h73;
		memory[16'h47f3] <= 8'h93;
		memory[16'h47f4] <= 8'h3a;
		memory[16'h47f5] <= 8'hcb;
		memory[16'h47f6] <= 8'h8e;
		memory[16'h47f7] <= 8'hf6;
		memory[16'h47f8] <= 8'h5;
		memory[16'h47f9] <= 8'h3d;
		memory[16'h47fa] <= 8'hee;
		memory[16'h47fb] <= 8'h61;
		memory[16'h47fc] <= 8'he4;
		memory[16'h47fd] <= 8'h5e;
		memory[16'h47fe] <= 8'h2c;
		memory[16'h47ff] <= 8'h5e;
		memory[16'h4800] <= 8'h1d;
		memory[16'h4801] <= 8'h12;
		memory[16'h4802] <= 8'h55;
		memory[16'h4803] <= 8'hf8;
		memory[16'h4804] <= 8'h80;
		memory[16'h4805] <= 8'hf8;
		memory[16'h4806] <= 8'hfe;
		memory[16'h4807] <= 8'hd8;
		memory[16'h4808] <= 8'h24;
		memory[16'h4809] <= 8'h45;
		memory[16'h480a] <= 8'h51;
		memory[16'h480b] <= 8'h2c;
		memory[16'h480c] <= 8'hb2;
		memory[16'h480d] <= 8'h40;
		memory[16'h480e] <= 8'h33;
		memory[16'h480f] <= 8'he1;
		memory[16'h4810] <= 8'h57;
		memory[16'h4811] <= 8'ha6;
		memory[16'h4812] <= 8'h74;
		memory[16'h4813] <= 8'h91;
		memory[16'h4814] <= 8'h72;
		memory[16'h4815] <= 8'h2;
		memory[16'h4816] <= 8'h87;
		memory[16'h4817] <= 8'h77;
		memory[16'h4818] <= 8'h40;
		memory[16'h4819] <= 8'h75;
		memory[16'h481a] <= 8'hd9;
		memory[16'h481b] <= 8'h24;
		memory[16'h481c] <= 8'hd4;
		memory[16'h481d] <= 8'h5;
		memory[16'h481e] <= 8'h83;
		memory[16'h481f] <= 8'hf1;
		memory[16'h4820] <= 8'h18;
		memory[16'h4821] <= 8'hd8;
		memory[16'h4822] <= 8'he9;
		memory[16'h4823] <= 8'h98;
		memory[16'h4824] <= 8'hd0;
		memory[16'h4825] <= 8'he7;
		memory[16'h4826] <= 8'h70;
		memory[16'h4827] <= 8'hf5;
		memory[16'h4828] <= 8'h2d;
		memory[16'h4829] <= 8'hc1;
		memory[16'h482a] <= 8'h21;
		memory[16'h482b] <= 8'hdf;
		memory[16'h482c] <= 8'h2;
		memory[16'h482d] <= 8'h54;
		memory[16'h482e] <= 8'hc0;
		memory[16'h482f] <= 8'h59;
		memory[16'h4830] <= 8'hfb;
		memory[16'h4831] <= 8'h34;
		memory[16'h4832] <= 8'hea;
		memory[16'h4833] <= 8'h6d;
		memory[16'h4834] <= 8'h37;
		memory[16'h4835] <= 8'h71;
		memory[16'h4836] <= 8'he4;
		memory[16'h4837] <= 8'h77;
		memory[16'h4838] <= 8'he7;
		memory[16'h4839] <= 8'hbd;
		memory[16'h483a] <= 8'h9b;
		memory[16'h483b] <= 8'hbb;
		memory[16'h483c] <= 8'hc3;
		memory[16'h483d] <= 8'h1e;
		memory[16'h483e] <= 8'hac;
		memory[16'h483f] <= 8'hdb;
		memory[16'h4840] <= 8'hf7;
		memory[16'h4841] <= 8'h95;
		memory[16'h4842] <= 8'h73;
		memory[16'h4843] <= 8'hc7;
		memory[16'h4844] <= 8'h7d;
		memory[16'h4845] <= 8'he4;
		memory[16'h4846] <= 8'hbc;
		memory[16'h4847] <= 8'haa;
		memory[16'h4848] <= 8'ha5;
		memory[16'h4849] <= 8'hde;
		memory[16'h484a] <= 8'h89;
		memory[16'h484b] <= 8'ha7;
		memory[16'h484c] <= 8'h32;
		memory[16'h484d] <= 8'h4a;
		memory[16'h484e] <= 8'h0;
		memory[16'h484f] <= 8'h2d;
		memory[16'h4850] <= 8'h7e;
		memory[16'h4851] <= 8'hea;
		memory[16'h4852] <= 8'h9a;
		memory[16'h4853] <= 8'hb5;
		memory[16'h4854] <= 8'h5c;
		memory[16'h4855] <= 8'h7f;
		memory[16'h4856] <= 8'h2c;
		memory[16'h4857] <= 8'h43;
		memory[16'h4858] <= 8'h3c;
		memory[16'h4859] <= 8'hc8;
		memory[16'h485a] <= 8'hfe;
		memory[16'h485b] <= 8'hff;
		memory[16'h485c] <= 8'he6;
		memory[16'h485d] <= 8'haa;
		memory[16'h485e] <= 8'hda;
		memory[16'h485f] <= 8'hdd;
		memory[16'h4860] <= 8'h3f;
		memory[16'h4861] <= 8'h4e;
		memory[16'h4862] <= 8'ha5;
		memory[16'h4863] <= 8'hbc;
		memory[16'h4864] <= 8'h32;
		memory[16'h4865] <= 8'h61;
		memory[16'h4866] <= 8'h66;
		memory[16'h4867] <= 8'hd7;
		memory[16'h4868] <= 8'h3f;
		memory[16'h4869] <= 8'hf0;
		memory[16'h486a] <= 8'h7f;
		memory[16'h486b] <= 8'h72;
		memory[16'h486c] <= 8'h3a;
		memory[16'h486d] <= 8'h7f;
		memory[16'h486e] <= 8'h9f;
		memory[16'h486f] <= 8'hb8;
		memory[16'h4870] <= 8'h6a;
		memory[16'h4871] <= 8'h3a;
		memory[16'h4872] <= 8'h6e;
		memory[16'h4873] <= 8'hc6;
		memory[16'h4874] <= 8'hb9;
		memory[16'h4875] <= 8'h9a;
		memory[16'h4876] <= 8'h9;
		memory[16'h4877] <= 8'hf5;
		memory[16'h4878] <= 8'h62;
		memory[16'h4879] <= 8'h7;
		memory[16'h487a] <= 8'hf5;
		memory[16'h487b] <= 8'h49;
		memory[16'h487c] <= 8'hb1;
		memory[16'h487d] <= 8'hcf;
		memory[16'h487e] <= 8'h26;
		memory[16'h487f] <= 8'hf0;
		memory[16'h4880] <= 8'h1d;
		memory[16'h4881] <= 8'hcb;
		memory[16'h4882] <= 8'had;
		memory[16'h4883] <= 8'h4f;
		memory[16'h4884] <= 8'h2d;
		memory[16'h4885] <= 8'h13;
		memory[16'h4886] <= 8'h27;
		memory[16'h4887] <= 8'h6c;
		memory[16'h4888] <= 8'h3;
		memory[16'h4889] <= 8'ha6;
		memory[16'h488a] <= 8'hde;
		memory[16'h488b] <= 8'h3d;
		memory[16'h488c] <= 8'h25;
		memory[16'h488d] <= 8'h7e;
		memory[16'h488e] <= 8'hf6;
		memory[16'h488f] <= 8'h8f;
		memory[16'h4890] <= 8'hb8;
		memory[16'h4891] <= 8'h64;
		memory[16'h4892] <= 8'h55;
		memory[16'h4893] <= 8'h71;
		memory[16'h4894] <= 8'hfe;
		memory[16'h4895] <= 8'h5e;
		memory[16'h4896] <= 8'h66;
		memory[16'h4897] <= 8'h61;
		memory[16'h4898] <= 8'h65;
		memory[16'h4899] <= 8'h5b;
		memory[16'h489a] <= 8'haa;
		memory[16'h489b] <= 8'h16;
		memory[16'h489c] <= 8'h2b;
		memory[16'h489d] <= 8'hd0;
		memory[16'h489e] <= 8'h7;
		memory[16'h489f] <= 8'h48;
		memory[16'h48a0] <= 8'h9c;
		memory[16'h48a1] <= 8'hb4;
		memory[16'h48a2] <= 8'h98;
		memory[16'h48a3] <= 8'hc9;
		memory[16'h48a4] <= 8'hc7;
		memory[16'h48a5] <= 8'hbf;
		memory[16'h48a6] <= 8'h35;
		memory[16'h48a7] <= 8'hcb;
		memory[16'h48a8] <= 8'h65;
		memory[16'h48a9] <= 8'h14;
		memory[16'h48aa] <= 8'h8;
		memory[16'h48ab] <= 8'h8a;
		memory[16'h48ac] <= 8'h92;
		memory[16'h48ad] <= 8'hfe;
		memory[16'h48ae] <= 8'h1a;
		memory[16'h48af] <= 8'h4a;
		memory[16'h48b0] <= 8'h62;
		memory[16'h48b1] <= 8'h6f;
		memory[16'h48b2] <= 8'hbb;
		memory[16'h48b3] <= 8'h61;
		memory[16'h48b4] <= 8'hce;
		memory[16'h48b5] <= 8'h21;
		memory[16'h48b6] <= 8'hc2;
		memory[16'h48b7] <= 8'h33;
		memory[16'h48b8] <= 8'h7d;
		memory[16'h48b9] <= 8'h6c;
		memory[16'h48ba] <= 8'h4a;
		memory[16'h48bb] <= 8'ha8;
		memory[16'h48bc] <= 8'h3c;
		memory[16'h48bd] <= 8'h51;
		memory[16'h48be] <= 8'hf0;
		memory[16'h48bf] <= 8'hd8;
		memory[16'h48c0] <= 8'h5;
		memory[16'h48c1] <= 8'h88;
		memory[16'h48c2] <= 8'ha1;
		memory[16'h48c3] <= 8'hcc;
		memory[16'h48c4] <= 8'h47;
		memory[16'h48c5] <= 8'hd7;
		memory[16'h48c6] <= 8'h97;
		memory[16'h48c7] <= 8'hac;
		memory[16'h48c8] <= 8'heb;
		memory[16'h48c9] <= 8'ha0;
		memory[16'h48ca] <= 8'h37;
		memory[16'h48cb] <= 8'h7d;
		memory[16'h48cc] <= 8'h9e;
		memory[16'h48cd] <= 8'h51;
		memory[16'h48ce] <= 8'hc7;
		memory[16'h48cf] <= 8'h1;
		memory[16'h48d0] <= 8'hc0;
		memory[16'h48d1] <= 8'h82;
		memory[16'h48d2] <= 8'h62;
		memory[16'h48d3] <= 8'h8e;
		memory[16'h48d4] <= 8'ha3;
		memory[16'h48d5] <= 8'h24;
		memory[16'h48d6] <= 8'hc2;
		memory[16'h48d7] <= 8'h20;
		memory[16'h48d8] <= 8'h90;
		memory[16'h48d9] <= 8'hc;
		memory[16'h48da] <= 8'hc8;
		memory[16'h48db] <= 8'hcc;
		memory[16'h48dc] <= 8'h5d;
		memory[16'h48dd] <= 8'hb9;
		memory[16'h48de] <= 8'ha5;
		memory[16'h48df] <= 8'h62;
		memory[16'h48e0] <= 8'h41;
		memory[16'h48e1] <= 8'h46;
		memory[16'h48e2] <= 8'h2e;
		memory[16'h48e3] <= 8'h89;
		memory[16'h48e4] <= 8'h1d;
		memory[16'h48e5] <= 8'hc6;
		memory[16'h48e6] <= 8'h35;
		memory[16'h48e7] <= 8'h8;
		memory[16'h48e8] <= 8'h66;
		memory[16'h48e9] <= 8'h6c;
		memory[16'h48ea] <= 8'h85;
		memory[16'h48eb] <= 8'h4;
		memory[16'h48ec] <= 8'hbd;
		memory[16'h48ed] <= 8'h4c;
		memory[16'h48ee] <= 8'h5;
		memory[16'h48ef] <= 8'h7e;
		memory[16'h48f0] <= 8'hce;
		memory[16'h48f1] <= 8'h67;
		memory[16'h48f2] <= 8'hc;
		memory[16'h48f3] <= 8'h72;
		memory[16'h48f4] <= 8'h8b;
		memory[16'h48f5] <= 8'hce;
		memory[16'h48f6] <= 8'h92;
		memory[16'h48f7] <= 8'h1b;
		memory[16'h48f8] <= 8'hda;
		memory[16'h48f9] <= 8'h5b;
		memory[16'h48fa] <= 8'he8;
		memory[16'h48fb] <= 8'h37;
		memory[16'h48fc] <= 8'h14;
		memory[16'h48fd] <= 8'h8d;
		memory[16'h48fe] <= 8'h99;
		memory[16'h48ff] <= 8'h55;
		memory[16'h4900] <= 8'hd3;
		memory[16'h4901] <= 8'hc8;
		memory[16'h4902] <= 8'hde;
		memory[16'h4903] <= 8'hf1;
		memory[16'h4904] <= 8'h8e;
		memory[16'h4905] <= 8'h14;
		memory[16'h4906] <= 8'hf9;
		memory[16'h4907] <= 8'hf4;
		memory[16'h4908] <= 8'h80;
		memory[16'h4909] <= 8'h7f;
		memory[16'h490a] <= 8'hf8;
		memory[16'h490b] <= 8'h3e;
		memory[16'h490c] <= 8'hcb;
		memory[16'h490d] <= 8'hfe;
		memory[16'h490e] <= 8'hbc;
		memory[16'h490f] <= 8'h9a;
		memory[16'h4910] <= 8'h65;
		memory[16'h4911] <= 8'hc8;
		memory[16'h4912] <= 8'hc;
		memory[16'h4913] <= 8'hf1;
		memory[16'h4914] <= 8'h97;
		memory[16'h4915] <= 8'h9e;
		memory[16'h4916] <= 8'hc;
		memory[16'h4917] <= 8'h71;
		memory[16'h4918] <= 8'hf9;
		memory[16'h4919] <= 8'hf4;
		memory[16'h491a] <= 8'ha9;
		memory[16'h491b] <= 8'hd;
		memory[16'h491c] <= 8'h81;
		memory[16'h491d] <= 8'h42;
		memory[16'h491e] <= 8'h63;
		memory[16'h491f] <= 8'h55;
		memory[16'h4920] <= 8'ha;
		memory[16'h4921] <= 8'h41;
		memory[16'h4922] <= 8'h46;
		memory[16'h4923] <= 8'h98;
		memory[16'h4924] <= 8'h55;
		memory[16'h4925] <= 8'h3f;
		memory[16'h4926] <= 8'h8c;
		memory[16'h4927] <= 8'hd6;
		memory[16'h4928] <= 8'hbe;
		memory[16'h4929] <= 8'h85;
		memory[16'h492a] <= 8'h14;
		memory[16'h492b] <= 8'h8a;
		memory[16'h492c] <= 8'h83;
		memory[16'h492d] <= 8'hd0;
		memory[16'h492e] <= 8'h24;
		memory[16'h492f] <= 8'he8;
		memory[16'h4930] <= 8'h98;
		memory[16'h4931] <= 8'h30;
		memory[16'h4932] <= 8'hd9;
		memory[16'h4933] <= 8'h2f;
		memory[16'h4934] <= 8'hce;
		memory[16'h4935] <= 8'he6;
		memory[16'h4936] <= 8'ha1;
		memory[16'h4937] <= 8'hc8;
		memory[16'h4938] <= 8'hda;
		memory[16'h4939] <= 8'h4a;
		memory[16'h493a] <= 8'hd5;
		memory[16'h493b] <= 8'h5c;
		memory[16'h493c] <= 8'h8c;
		memory[16'h493d] <= 8'h38;
		memory[16'h493e] <= 8'hb1;
		memory[16'h493f] <= 8'h97;
		memory[16'h4940] <= 8'h7a;
		memory[16'h4941] <= 8'hf7;
		memory[16'h4942] <= 8'h2f;
		memory[16'h4943] <= 8'hcf;
		memory[16'h4944] <= 8'h36;
		memory[16'h4945] <= 8'hbc;
		memory[16'h4946] <= 8'ha5;
		memory[16'h4947] <= 8'hf5;
		memory[16'h4948] <= 8'h41;
		memory[16'h4949] <= 8'hb9;
		memory[16'h494a] <= 8'h7f;
		memory[16'h494b] <= 8'hc4;
		memory[16'h494c] <= 8'h89;
		memory[16'h494d] <= 8'ha3;
		memory[16'h494e] <= 8'hac;
		memory[16'h494f] <= 8'h22;
		memory[16'h4950] <= 8'hd3;
		memory[16'h4951] <= 8'h86;
		memory[16'h4952] <= 8'h51;
		memory[16'h4953] <= 8'ha1;
		memory[16'h4954] <= 8'h6c;
		memory[16'h4955] <= 8'hf2;
		memory[16'h4956] <= 8'h69;
		memory[16'h4957] <= 8'h46;
		memory[16'h4958] <= 8'h3c;
		memory[16'h4959] <= 8'h3f;
		memory[16'h495a] <= 8'ha2;
		memory[16'h495b] <= 8'hc9;
		memory[16'h495c] <= 8'h77;
		memory[16'h495d] <= 8'h53;
		memory[16'h495e] <= 8'h60;
		memory[16'h495f] <= 8'hf1;
		memory[16'h4960] <= 8'h4a;
		memory[16'h4961] <= 8'h8f;
		memory[16'h4962] <= 8'hc1;
		memory[16'h4963] <= 8'h81;
		memory[16'h4964] <= 8'h4b;
		memory[16'h4965] <= 8'h66;
		memory[16'h4966] <= 8'h76;
		memory[16'h4967] <= 8'h8c;
		memory[16'h4968] <= 8'h20;
		memory[16'h4969] <= 8'hf5;
		memory[16'h496a] <= 8'h50;
		memory[16'h496b] <= 8'ha9;
		memory[16'h496c] <= 8'h98;
		memory[16'h496d] <= 8'hfd;
		memory[16'h496e] <= 8'hcb;
		memory[16'h496f] <= 8'h6b;
		memory[16'h4970] <= 8'h83;
		memory[16'h4971] <= 8'h1d;
		memory[16'h4972] <= 8'hc;
		memory[16'h4973] <= 8'hef;
		memory[16'h4974] <= 8'hf;
		memory[16'h4975] <= 8'h76;
		memory[16'h4976] <= 8'h35;
		memory[16'h4977] <= 8'h4c;
		memory[16'h4978] <= 8'hb5;
		memory[16'h4979] <= 8'hd8;
		memory[16'h497a] <= 8'h15;
		memory[16'h497b] <= 8'h2c;
		memory[16'h497c] <= 8'h2b;
		memory[16'h497d] <= 8'h75;
		memory[16'h497e] <= 8'h1e;
		memory[16'h497f] <= 8'h76;
		memory[16'h4980] <= 8'h4;
		memory[16'h4981] <= 8'hdf;
		memory[16'h4982] <= 8'hf7;
		memory[16'h4983] <= 8'h50;
		memory[16'h4984] <= 8'h45;
		memory[16'h4985] <= 8'h6d;
		memory[16'h4986] <= 8'hdc;
		memory[16'h4987] <= 8'h65;
		memory[16'h4988] <= 8'h62;
		memory[16'h4989] <= 8'h2d;
		memory[16'h498a] <= 8'hf;
		memory[16'h498b] <= 8'hfa;
		memory[16'h498c] <= 8'h2a;
		memory[16'h498d] <= 8'hda;
		memory[16'h498e] <= 8'h65;
		memory[16'h498f] <= 8'had;
		memory[16'h4990] <= 8'hf7;
		memory[16'h4991] <= 8'h71;
		memory[16'h4992] <= 8'h9c;
		memory[16'h4993] <= 8'h7;
		memory[16'h4994] <= 8'he7;
		memory[16'h4995] <= 8'hd1;
		memory[16'h4996] <= 8'h53;
		memory[16'h4997] <= 8'h9c;
		memory[16'h4998] <= 8'ha9;
		memory[16'h4999] <= 8'h68;
		memory[16'h499a] <= 8'hc9;
		memory[16'h499b] <= 8'hd5;
		memory[16'h499c] <= 8'hdd;
		memory[16'h499d] <= 8'he7;
		memory[16'h499e] <= 8'h4b;
		memory[16'h499f] <= 8'he1;
		memory[16'h49a0] <= 8'hc6;
		memory[16'h49a1] <= 8'h42;
		memory[16'h49a2] <= 8'h31;
		memory[16'h49a3] <= 8'hb;
		memory[16'h49a4] <= 8'haf;
		memory[16'h49a5] <= 8'he;
		memory[16'h49a6] <= 8'h71;
		memory[16'h49a7] <= 8'h11;
		memory[16'h49a8] <= 8'h3b;
		memory[16'h49a9] <= 8'h80;
		memory[16'h49aa] <= 8'hb;
		memory[16'h49ab] <= 8'h65;
		memory[16'h49ac] <= 8'h5a;
		memory[16'h49ad] <= 8'h70;
		memory[16'h49ae] <= 8'h12;
		memory[16'h49af] <= 8'h52;
		memory[16'h49b0] <= 8'he1;
		memory[16'h49b1] <= 8'hae;
		memory[16'h49b2] <= 8'h59;
		memory[16'h49b3] <= 8'hc9;
		memory[16'h49b4] <= 8'h7f;
		memory[16'h49b5] <= 8'hac;
		memory[16'h49b6] <= 8'h65;
		memory[16'h49b7] <= 8'h29;
		memory[16'h49b8] <= 8'h14;
		memory[16'h49b9] <= 8'h2e;
		memory[16'h49ba] <= 8'hfe;
		memory[16'h49bb] <= 8'hf1;
		memory[16'h49bc] <= 8'h15;
		memory[16'h49bd] <= 8'h49;
		memory[16'h49be] <= 8'hd2;
		memory[16'h49bf] <= 8'hdb;
		memory[16'h49c0] <= 8'h8b;
		memory[16'h49c1] <= 8'h4;
		memory[16'h49c2] <= 8'he7;
		memory[16'h49c3] <= 8'h3a;
		memory[16'h49c4] <= 8'h12;
		memory[16'h49c5] <= 8'h58;
		memory[16'h49c6] <= 8'h4b;
		memory[16'h49c7] <= 8'h4d;
		memory[16'h49c8] <= 8'hd8;
		memory[16'h49c9] <= 8'h56;
		memory[16'h49ca] <= 8'hb2;
		memory[16'h49cb] <= 8'h32;
		memory[16'h49cc] <= 8'hc6;
		memory[16'h49cd] <= 8'hc4;
		memory[16'h49ce] <= 8'h84;
		memory[16'h49cf] <= 8'ha7;
		memory[16'h49d0] <= 8'h72;
		memory[16'h49d1] <= 8'hdd;
		memory[16'h49d2] <= 8'h70;
		memory[16'h49d3] <= 8'hf1;
		memory[16'h49d4] <= 8'h89;
		memory[16'h49d5] <= 8'hd6;
		memory[16'h49d6] <= 8'h1a;
		memory[16'h49d7] <= 8'h9d;
		memory[16'h49d8] <= 8'h4;
		memory[16'h49d9] <= 8'h18;
		memory[16'h49da] <= 8'h8e;
		memory[16'h49db] <= 8'h1a;
		memory[16'h49dc] <= 8'h61;
		memory[16'h49dd] <= 8'h61;
		memory[16'h49de] <= 8'hf5;
		memory[16'h49df] <= 8'hec;
		memory[16'h49e0] <= 8'h65;
		memory[16'h49e1] <= 8'hdc;
		memory[16'h49e2] <= 8'h26;
		memory[16'h49e3] <= 8'h77;
		memory[16'h49e4] <= 8'h34;
		memory[16'h49e5] <= 8'h71;
		memory[16'h49e6] <= 8'hc4;
		memory[16'h49e7] <= 8'hc;
		memory[16'h49e8] <= 8'hc7;
		memory[16'h49e9] <= 8'h76;
		memory[16'h49ea] <= 8'h3f;
		memory[16'h49eb] <= 8'h8d;
		memory[16'h49ec] <= 8'h3a;
		memory[16'h49ed] <= 8'hc3;
		memory[16'h49ee] <= 8'h35;
		memory[16'h49ef] <= 8'hac;
		memory[16'h49f0] <= 8'ha1;
		memory[16'h49f1] <= 8'ha5;
		memory[16'h49f2] <= 8'h9d;
		memory[16'h49f3] <= 8'h2a;
		memory[16'h49f4] <= 8'h7b;
		memory[16'h49f5] <= 8'hb8;
		memory[16'h49f6] <= 8'hc8;
		memory[16'h49f7] <= 8'h80;
		memory[16'h49f8] <= 8'hd0;
		memory[16'h49f9] <= 8'h56;
		memory[16'h49fa] <= 8'h9a;
		memory[16'h49fb] <= 8'h32;
		memory[16'h49fc] <= 8'hb7;
		memory[16'h49fd] <= 8'h8f;
		memory[16'h49fe] <= 8'h1e;
		memory[16'h49ff] <= 8'h1c;
		memory[16'h4a00] <= 8'h6c;
		memory[16'h4a01] <= 8'h45;
		memory[16'h4a02] <= 8'h93;
		memory[16'h4a03] <= 8'ha0;
		memory[16'h4a04] <= 8'hb6;
		memory[16'h4a05] <= 8'h57;
		memory[16'h4a06] <= 8'had;
		memory[16'h4a07] <= 8'h7e;
		memory[16'h4a08] <= 8'hcd;
		memory[16'h4a09] <= 8'hec;
		memory[16'h4a0a] <= 8'hb;
		memory[16'h4a0b] <= 8'h7;
		memory[16'h4a0c] <= 8'haf;
		memory[16'h4a0d] <= 8'h40;
		memory[16'h4a0e] <= 8'hb3;
		memory[16'h4a0f] <= 8'h50;
		memory[16'h4a10] <= 8'he6;
		memory[16'h4a11] <= 8'h51;
		memory[16'h4a12] <= 8'h7b;
		memory[16'h4a13] <= 8'h61;
		memory[16'h4a14] <= 8'h9;
		memory[16'h4a15] <= 8'h43;
		memory[16'h4a16] <= 8'he1;
		memory[16'h4a17] <= 8'hd9;
		memory[16'h4a18] <= 8'h99;
		memory[16'h4a19] <= 8'h7b;
		memory[16'h4a1a] <= 8'hb;
		memory[16'h4a1b] <= 8'h51;
		memory[16'h4a1c] <= 8'hb;
		memory[16'h4a1d] <= 8'h2a;
		memory[16'h4a1e] <= 8'h6d;
		memory[16'h4a1f] <= 8'h77;
		memory[16'h4a20] <= 8'h6f;
		memory[16'h4a21] <= 8'h1;
		memory[16'h4a22] <= 8'h17;
		memory[16'h4a23] <= 8'h25;
		memory[16'h4a24] <= 8'h58;
		memory[16'h4a25] <= 8'hc4;
		memory[16'h4a26] <= 8'ha3;
		memory[16'h4a27] <= 8'h26;
		memory[16'h4a28] <= 8'hb0;
		memory[16'h4a29] <= 8'haf;
		memory[16'h4a2a] <= 8'h2d;
		memory[16'h4a2b] <= 8'h60;
		memory[16'h4a2c] <= 8'hef;
		memory[16'h4a2d] <= 8'he1;
		memory[16'h4a2e] <= 8'hb0;
		memory[16'h4a2f] <= 8'hd5;
		memory[16'h4a30] <= 8'h32;
		memory[16'h4a31] <= 8'h2b;
		memory[16'h4a32] <= 8'h37;
		memory[16'h4a33] <= 8'h3b;
		memory[16'h4a34] <= 8'h6e;
		memory[16'h4a35] <= 8'h18;
		memory[16'h4a36] <= 8'h14;
		memory[16'h4a37] <= 8'h8;
		memory[16'h4a38] <= 8'h94;
		memory[16'h4a39] <= 8'h20;
		memory[16'h4a3a] <= 8'h59;
		memory[16'h4a3b] <= 8'h9f;
		memory[16'h4a3c] <= 8'h4a;
		memory[16'h4a3d] <= 8'hc6;
		memory[16'h4a3e] <= 8'h16;
		memory[16'h4a3f] <= 8'hb9;
		memory[16'h4a40] <= 8'hc7;
		memory[16'h4a41] <= 8'h2d;
		memory[16'h4a42] <= 8'hde;
		memory[16'h4a43] <= 8'h20;
		memory[16'h4a44] <= 8'hf2;
		memory[16'h4a45] <= 8'h82;
		memory[16'h4a46] <= 8'h46;
		memory[16'h4a47] <= 8'ha2;
		memory[16'h4a48] <= 8'h31;
		memory[16'h4a49] <= 8'h73;
		memory[16'h4a4a] <= 8'h2;
		memory[16'h4a4b] <= 8'h20;
		memory[16'h4a4c] <= 8'h54;
		memory[16'h4a4d] <= 8'hb3;
		memory[16'h4a4e] <= 8'hf6;
		memory[16'h4a4f] <= 8'h86;
		memory[16'h4a50] <= 8'hde;
		memory[16'h4a51] <= 8'h2d;
		memory[16'h4a52] <= 8'hc1;
		memory[16'h4a53] <= 8'h4d;
		memory[16'h4a54] <= 8'h45;
		memory[16'h4a55] <= 8'hd6;
		memory[16'h4a56] <= 8'h55;
		memory[16'h4a57] <= 8'hd9;
		memory[16'h4a58] <= 8'hf6;
		memory[16'h4a59] <= 8'hae;
		memory[16'h4a5a] <= 8'h78;
		memory[16'h4a5b] <= 8'h40;
		memory[16'h4a5c] <= 8'h74;
		memory[16'h4a5d] <= 8'h8e;
		memory[16'h4a5e] <= 8'hf9;
		memory[16'h4a5f] <= 8'h3c;
		memory[16'h4a60] <= 8'hbc;
		memory[16'h4a61] <= 8'hd7;
		memory[16'h4a62] <= 8'h5c;
		memory[16'h4a63] <= 8'hae;
		memory[16'h4a64] <= 8'h59;
		memory[16'h4a65] <= 8'ha2;
		memory[16'h4a66] <= 8'h50;
		memory[16'h4a67] <= 8'h8a;
		memory[16'h4a68] <= 8'h15;
		memory[16'h4a69] <= 8'h53;
		memory[16'h4a6a] <= 8'hab;
		memory[16'h4a6b] <= 8'h6a;
		memory[16'h4a6c] <= 8'h6;
		memory[16'h4a6d] <= 8'ha1;
		memory[16'h4a6e] <= 8'hf0;
		memory[16'h4a6f] <= 8'he4;
		memory[16'h4a70] <= 8'hce;
		memory[16'h4a71] <= 8'hb2;
		memory[16'h4a72] <= 8'h31;
		memory[16'h4a73] <= 8'h13;
		memory[16'h4a74] <= 8'h88;
		memory[16'h4a75] <= 8'h86;
		memory[16'h4a76] <= 8'hed;
		memory[16'h4a77] <= 8'h7e;
		memory[16'h4a78] <= 8'h34;
		memory[16'h4a79] <= 8'h65;
		memory[16'h4a7a] <= 8'hbe;
		memory[16'h4a7b] <= 8'ha9;
		memory[16'h4a7c] <= 8'hf4;
		memory[16'h4a7d] <= 8'hb7;
		memory[16'h4a7e] <= 8'he5;
		memory[16'h4a7f] <= 8'hb0;
		memory[16'h4a80] <= 8'h8e;
		memory[16'h4a81] <= 8'h41;
		memory[16'h4a82] <= 8'h5e;
		memory[16'h4a83] <= 8'he8;
		memory[16'h4a84] <= 8'he3;
		memory[16'h4a85] <= 8'hae;
		memory[16'h4a86] <= 8'h72;
		memory[16'h4a87] <= 8'hf8;
		memory[16'h4a88] <= 8'h1;
		memory[16'h4a89] <= 8'h1d;
		memory[16'h4a8a] <= 8'h62;
		memory[16'h4a8b] <= 8'h7;
		memory[16'h4a8c] <= 8'hbe;
		memory[16'h4a8d] <= 8'h53;
		memory[16'h4a8e] <= 8'hec;
		memory[16'h4a8f] <= 8'h8c;
		memory[16'h4a90] <= 8'h5;
		memory[16'h4a91] <= 8'h1d;
		memory[16'h4a92] <= 8'ha0;
		memory[16'h4a93] <= 8'h8d;
		memory[16'h4a94] <= 8'ha4;
		memory[16'h4a95] <= 8'h8d;
		memory[16'h4a96] <= 8'hb;
		memory[16'h4a97] <= 8'hd8;
		memory[16'h4a98] <= 8'hf2;
		memory[16'h4a99] <= 8'hc9;
		memory[16'h4a9a] <= 8'h81;
		memory[16'h4a9b] <= 8'he6;
		memory[16'h4a9c] <= 8'h80;
		memory[16'h4a9d] <= 8'h66;
		memory[16'h4a9e] <= 8'h96;
		memory[16'h4a9f] <= 8'he;
		memory[16'h4aa0] <= 8'ha7;
		memory[16'h4aa1] <= 8'hf4;
		memory[16'h4aa2] <= 8'hf6;
		memory[16'h4aa3] <= 8'h8a;
		memory[16'h4aa4] <= 8'ha3;
		memory[16'h4aa5] <= 8'h69;
		memory[16'h4aa6] <= 8'h83;
		memory[16'h4aa7] <= 8'ha4;
		memory[16'h4aa8] <= 8'h86;
		memory[16'h4aa9] <= 8'he5;
		memory[16'h4aaa] <= 8'hac;
		memory[16'h4aab] <= 8'h45;
		memory[16'h4aac] <= 8'h38;
		memory[16'h4aad] <= 8'h98;
		memory[16'h4aae] <= 8'hd1;
		memory[16'h4aaf] <= 8'h3d;
		memory[16'h4ab0] <= 8'hb5;
		memory[16'h4ab1] <= 8'h71;
		memory[16'h4ab2] <= 8'hca;
		memory[16'h4ab3] <= 8'h59;
		memory[16'h4ab4] <= 8'hfe;
		memory[16'h4ab5] <= 8'hd5;
		memory[16'h4ab6] <= 8'h32;
		memory[16'h4ab7] <= 8'hf1;
		memory[16'h4ab8] <= 8'h9e;
		memory[16'h4ab9] <= 8'hb3;
		memory[16'h4aba] <= 8'hd7;
		memory[16'h4abb] <= 8'h1e;
		memory[16'h4abc] <= 8'h1a;
		memory[16'h4abd] <= 8'h6e;
		memory[16'h4abe] <= 8'h2d;
		memory[16'h4abf] <= 8'hc1;
		memory[16'h4ac0] <= 8'h62;
		memory[16'h4ac1] <= 8'h23;
		memory[16'h4ac2] <= 8'h4c;
		memory[16'h4ac3] <= 8'h5;
		memory[16'h4ac4] <= 8'h8c;
		memory[16'h4ac5] <= 8'hcf;
		memory[16'h4ac6] <= 8'haa;
		memory[16'h4ac7] <= 8'h13;
		memory[16'h4ac8] <= 8'hb4;
		memory[16'h4ac9] <= 8'h56;
		memory[16'h4aca] <= 8'h58;
		memory[16'h4acb] <= 8'hed;
		memory[16'h4acc] <= 8'hee;
		memory[16'h4acd] <= 8'h29;
		memory[16'h4ace] <= 8'h2a;
		memory[16'h4acf] <= 8'ha3;
		memory[16'h4ad0] <= 8'h9b;
		memory[16'h4ad1] <= 8'hf5;
		memory[16'h4ad2] <= 8'hfd;
		memory[16'h4ad3] <= 8'h99;
		memory[16'h4ad4] <= 8'hca;
		memory[16'h4ad5] <= 8'h2f;
		memory[16'h4ad6] <= 8'h8a;
		memory[16'h4ad7] <= 8'h69;
		memory[16'h4ad8] <= 8'he2;
		memory[16'h4ad9] <= 8'h62;
		memory[16'h4ada] <= 8'h87;
		memory[16'h4adb] <= 8'hfc;
		memory[16'h4adc] <= 8'hd0;
		memory[16'h4add] <= 8'hb4;
		memory[16'h4ade] <= 8'hbe;
		memory[16'h4adf] <= 8'h32;
		memory[16'h4ae0] <= 8'hd8;
		memory[16'h4ae1] <= 8'ha;
		memory[16'h4ae2] <= 8'h38;
		memory[16'h4ae3] <= 8'h64;
		memory[16'h4ae4] <= 8'hd9;
		memory[16'h4ae5] <= 8'he2;
		memory[16'h4ae6] <= 8'h77;
		memory[16'h4ae7] <= 8'h8d;
		memory[16'h4ae8] <= 8'h38;
		memory[16'h4ae9] <= 8'hcf;
		memory[16'h4aea] <= 8'h7a;
		memory[16'h4aeb] <= 8'h26;
		memory[16'h4aec] <= 8'hf9;
		memory[16'h4aed] <= 8'ha5;
		memory[16'h4aee] <= 8'hc9;
		memory[16'h4aef] <= 8'h94;
		memory[16'h4af0] <= 8'h9a;
		memory[16'h4af1] <= 8'hc6;
		memory[16'h4af2] <= 8'h2d;
		memory[16'h4af3] <= 8'h64;
		memory[16'h4af4] <= 8'hf5;
		memory[16'h4af5] <= 8'hb8;
		memory[16'h4af6] <= 8'hcd;
		memory[16'h4af7] <= 8'hd8;
		memory[16'h4af8] <= 8'h1a;
		memory[16'h4af9] <= 8'h55;
		memory[16'h4afa] <= 8'hd4;
		memory[16'h4afb] <= 8'hea;
		memory[16'h4afc] <= 8'h9;
		memory[16'h4afd] <= 8'h92;
		memory[16'h4afe] <= 8'h1c;
		memory[16'h4aff] <= 8'he1;
		memory[16'h4b00] <= 8'h9c;
		memory[16'h4b01] <= 8'h54;
		memory[16'h4b02] <= 8'h46;
		memory[16'h4b03] <= 8'h75;
		memory[16'h4b04] <= 8'h36;
		memory[16'h4b05] <= 8'hbd;
		memory[16'h4b06] <= 8'h3;
		memory[16'h4b07] <= 8'h6e;
		memory[16'h4b08] <= 8'h8d;
		memory[16'h4b09] <= 8'h7d;
		memory[16'h4b0a] <= 8'h94;
		memory[16'h4b0b] <= 8'h86;
		memory[16'h4b0c] <= 8'h22;
		memory[16'h4b0d] <= 8'h5e;
		memory[16'h4b0e] <= 8'h1a;
		memory[16'h4b0f] <= 8'hbc;
		memory[16'h4b10] <= 8'h24;
		memory[16'h4b11] <= 8'h47;
		memory[16'h4b12] <= 8'h21;
		memory[16'h4b13] <= 8'h1a;
		memory[16'h4b14] <= 8'hff;
		memory[16'h4b15] <= 8'hee;
		memory[16'h4b16] <= 8'hf2;
		memory[16'h4b17] <= 8'h19;
		memory[16'h4b18] <= 8'h43;
		memory[16'h4b19] <= 8'hc6;
		memory[16'h4b1a] <= 8'h3;
		memory[16'h4b1b] <= 8'h4d;
		memory[16'h4b1c] <= 8'h59;
		memory[16'h4b1d] <= 8'h20;
		memory[16'h4b1e] <= 8'h2e;
		memory[16'h4b1f] <= 8'hf5;
		memory[16'h4b20] <= 8'h74;
		memory[16'h4b21] <= 8'h74;
		memory[16'h4b22] <= 8'h6b;
		memory[16'h4b23] <= 8'hab;
		memory[16'h4b24] <= 8'h32;
		memory[16'h4b25] <= 8'h6e;
		memory[16'h4b26] <= 8'h19;
		memory[16'h4b27] <= 8'hbf;
		memory[16'h4b28] <= 8'heb;
		memory[16'h4b29] <= 8'hae;
		memory[16'h4b2a] <= 8'h45;
		memory[16'h4b2b] <= 8'he;
		memory[16'h4b2c] <= 8'hc;
		memory[16'h4b2d] <= 8'h5f;
		memory[16'h4b2e] <= 8'hca;
		memory[16'h4b2f] <= 8'h30;
		memory[16'h4b30] <= 8'ha6;
		memory[16'h4b31] <= 8'heb;
		memory[16'h4b32] <= 8'h4a;
		memory[16'h4b33] <= 8'ha6;
		memory[16'h4b34] <= 8'hda;
		memory[16'h4b35] <= 8'h3c;
		memory[16'h4b36] <= 8'hbf;
		memory[16'h4b37] <= 8'h1d;
		memory[16'h4b38] <= 8'h3;
		memory[16'h4b39] <= 8'hc3;
		memory[16'h4b3a] <= 8'h6a;
		memory[16'h4b3b] <= 8'h5c;
		memory[16'h4b3c] <= 8'he3;
		memory[16'h4b3d] <= 8'h99;
		memory[16'h4b3e] <= 8'h51;
		memory[16'h4b3f] <= 8'h57;
		memory[16'h4b40] <= 8'hd;
		memory[16'h4b41] <= 8'hbc;
		memory[16'h4b42] <= 8'h2;
		memory[16'h4b43] <= 8'h3f;
		memory[16'h4b44] <= 8'h2a;
		memory[16'h4b45] <= 8'h1c;
		memory[16'h4b46] <= 8'hfe;
		memory[16'h4b47] <= 8'h16;
		memory[16'h4b48] <= 8'hca;
		memory[16'h4b49] <= 8'h43;
		memory[16'h4b4a] <= 8'h24;
		memory[16'h4b4b] <= 8'hd6;
		memory[16'h4b4c] <= 8'ha2;
		memory[16'h4b4d] <= 8'hee;
		memory[16'h4b4e] <= 8'h6;
		memory[16'h4b4f] <= 8'h49;
		memory[16'h4b50] <= 8'hda;
		memory[16'h4b51] <= 8'h51;
		memory[16'h4b52] <= 8'hef;
		memory[16'h4b53] <= 8'hb4;
		memory[16'h4b54] <= 8'h8d;
		memory[16'h4b55] <= 8'hae;
		memory[16'h4b56] <= 8'hd1;
		memory[16'h4b57] <= 8'h90;
		memory[16'h4b58] <= 8'h71;
		memory[16'h4b59] <= 8'h3c;
		memory[16'h4b5a] <= 8'hec;
		memory[16'h4b5b] <= 8'h54;
		memory[16'h4b5c] <= 8'hd5;
		memory[16'h4b5d] <= 8'h3e;
		memory[16'h4b5e] <= 8'hac;
		memory[16'h4b5f] <= 8'he2;
		memory[16'h4b60] <= 8'hfa;
		memory[16'h4b61] <= 8'hae;
		memory[16'h4b62] <= 8'h22;
		memory[16'h4b63] <= 8'h25;
		memory[16'h4b64] <= 8'hca;
		memory[16'h4b65] <= 8'h20;
		memory[16'h4b66] <= 8'h3b;
		memory[16'h4b67] <= 8'h94;
		memory[16'h4b68] <= 8'h64;
		memory[16'h4b69] <= 8'h5f;
		memory[16'h4b6a] <= 8'h6a;
		memory[16'h4b6b] <= 8'h6;
		memory[16'h4b6c] <= 8'h4d;
		memory[16'h4b6d] <= 8'h71;
		memory[16'h4b6e] <= 8'h4f;
		memory[16'h4b6f] <= 8'h27;
		memory[16'h4b70] <= 8'hc2;
		memory[16'h4b71] <= 8'h3e;
		memory[16'h4b72] <= 8'hdb;
		memory[16'h4b73] <= 8'h4f;
		memory[16'h4b74] <= 8'hed;
		memory[16'h4b75] <= 8'had;
		memory[16'h4b76] <= 8'he0;
		memory[16'h4b77] <= 8'h5e;
		memory[16'h4b78] <= 8'he9;
		memory[16'h4b79] <= 8'hcc;
		memory[16'h4b7a] <= 8'hb3;
		memory[16'h4b7b] <= 8'hbe;
		memory[16'h4b7c] <= 8'ha;
		memory[16'h4b7d] <= 8'h5f;
		memory[16'h4b7e] <= 8'ha0;
		memory[16'h4b7f] <= 8'h5;
		memory[16'h4b80] <= 8'hd;
		memory[16'h4b81] <= 8'hc2;
		memory[16'h4b82] <= 8'h2a;
		memory[16'h4b83] <= 8'hd8;
		memory[16'h4b84] <= 8'he3;
		memory[16'h4b85] <= 8'h65;
		memory[16'h4b86] <= 8'h6c;
		memory[16'h4b87] <= 8'h47;
		memory[16'h4b88] <= 8'hc4;
		memory[16'h4b89] <= 8'hd7;
		memory[16'h4b8a] <= 8'h4d;
		memory[16'h4b8b] <= 8'h11;
		memory[16'h4b8c] <= 8'h48;
		memory[16'h4b8d] <= 8'h9d;
		memory[16'h4b8e] <= 8'h39;
		memory[16'h4b8f] <= 8'ha;
		memory[16'h4b90] <= 8'hdb;
		memory[16'h4b91] <= 8'h14;
		memory[16'h4b92] <= 8'h59;
		memory[16'h4b93] <= 8'hc8;
		memory[16'h4b94] <= 8'hc1;
		memory[16'h4b95] <= 8'h39;
		memory[16'h4b96] <= 8'h27;
		memory[16'h4b97] <= 8'haa;
		memory[16'h4b98] <= 8'h6;
		memory[16'h4b99] <= 8'hda;
		memory[16'h4b9a] <= 8'h68;
		memory[16'h4b9b] <= 8'h10;
		memory[16'h4b9c] <= 8'h39;
		memory[16'h4b9d] <= 8'h9;
		memory[16'h4b9e] <= 8'h15;
		memory[16'h4b9f] <= 8'h46;
		memory[16'h4ba0] <= 8'hcb;
		memory[16'h4ba1] <= 8'h3f;
		memory[16'h4ba2] <= 8'h1e;
		memory[16'h4ba3] <= 8'hae;
		memory[16'h4ba4] <= 8'ha4;
		memory[16'h4ba5] <= 8'h8b;
		memory[16'h4ba6] <= 8'hf5;
		memory[16'h4ba7] <= 8'h68;
		memory[16'h4ba8] <= 8'h62;
		memory[16'h4ba9] <= 8'h43;
		memory[16'h4baa] <= 8'h7a;
		memory[16'h4bab] <= 8'haa;
		memory[16'h4bac] <= 8'he0;
		memory[16'h4bad] <= 8'hb3;
		memory[16'h4bae] <= 8'hb4;
		memory[16'h4baf] <= 8'hbb;
		memory[16'h4bb0] <= 8'hc7;
		memory[16'h4bb1] <= 8'hd;
		memory[16'h4bb2] <= 8'h84;
		memory[16'h4bb3] <= 8'h89;
		memory[16'h4bb4] <= 8'h47;
		memory[16'h4bb5] <= 8'hab;
		memory[16'h4bb6] <= 8'h33;
		memory[16'h4bb7] <= 8'h4d;
		memory[16'h4bb8] <= 8'h85;
		memory[16'h4bb9] <= 8'h9c;
		memory[16'h4bba] <= 8'h5d;
		memory[16'h4bbb] <= 8'hbe;
		memory[16'h4bbc] <= 8'ha5;
		memory[16'h4bbd] <= 8'h73;
		memory[16'h4bbe] <= 8'h4;
		memory[16'h4bbf] <= 8'h70;
		memory[16'h4bc0] <= 8'hb2;
		memory[16'h4bc1] <= 8'h23;
		memory[16'h4bc2] <= 8'h1f;
		memory[16'h4bc3] <= 8'h57;
		memory[16'h4bc4] <= 8'hae;
		memory[16'h4bc5] <= 8'h14;
		memory[16'h4bc6] <= 8'hbf;
		memory[16'h4bc7] <= 8'h10;
		memory[16'h4bc8] <= 8'h57;
		memory[16'h4bc9] <= 8'h39;
		memory[16'h4bca] <= 8'hba;
		memory[16'h4bcb] <= 8'h37;
		memory[16'h4bcc] <= 8'hec;
		memory[16'h4bcd] <= 8'h6e;
		memory[16'h4bce] <= 8'hf3;
		memory[16'h4bcf] <= 8'hb4;
		memory[16'h4bd0] <= 8'h7b;
		memory[16'h4bd1] <= 8'h77;
		memory[16'h4bd2] <= 8'h3d;
		memory[16'h4bd3] <= 8'hc2;
		memory[16'h4bd4] <= 8'h22;
		memory[16'h4bd5] <= 8'h70;
		memory[16'h4bd6] <= 8'hf;
		memory[16'h4bd7] <= 8'ha7;
		memory[16'h4bd8] <= 8'hc;
		memory[16'h4bd9] <= 8'h6d;
		memory[16'h4bda] <= 8'h65;
		memory[16'h4bdb] <= 8'hb1;
		memory[16'h4bdc] <= 8'he0;
		memory[16'h4bdd] <= 8'h69;
		memory[16'h4bde] <= 8'h22;
		memory[16'h4bdf] <= 8'h92;
		memory[16'h4be0] <= 8'h8c;
		memory[16'h4be1] <= 8'h41;
		memory[16'h4be2] <= 8'he9;
		memory[16'h4be3] <= 8'h3a;
		memory[16'h4be4] <= 8'h55;
		memory[16'h4be5] <= 8'ha9;
		memory[16'h4be6] <= 8'h4a;
		memory[16'h4be7] <= 8'had;
		memory[16'h4be8] <= 8'he2;
		memory[16'h4be9] <= 8'h4;
		memory[16'h4bea] <= 8'he4;
		memory[16'h4beb] <= 8'hcf;
		memory[16'h4bec] <= 8'h72;
		memory[16'h4bed] <= 8'hd7;
		memory[16'h4bee] <= 8'h83;
		memory[16'h4bef] <= 8'hee;
		memory[16'h4bf0] <= 8'h4e;
		memory[16'h4bf1] <= 8'hc0;
		memory[16'h4bf2] <= 8'hb0;
		memory[16'h4bf3] <= 8'h70;
		memory[16'h4bf4] <= 8'h30;
		memory[16'h4bf5] <= 8'hc0;
		memory[16'h4bf6] <= 8'h17;
		memory[16'h4bf7] <= 8'h3d;
		memory[16'h4bf8] <= 8'h2d;
		memory[16'h4bf9] <= 8'h7c;
		memory[16'h4bfa] <= 8'hee;
		memory[16'h4bfb] <= 8'hd;
		memory[16'h4bfc] <= 8'he6;
		memory[16'h4bfd] <= 8'h10;
		memory[16'h4bfe] <= 8'h9f;
		memory[16'h4bff] <= 8'h72;
		memory[16'h4c00] <= 8'h51;
		memory[16'h4c01] <= 8'h89;
		memory[16'h4c02] <= 8'had;
		memory[16'h4c03] <= 8'ha7;
		memory[16'h4c04] <= 8'h32;
		memory[16'h4c05] <= 8'hf7;
		memory[16'h4c06] <= 8'h54;
		memory[16'h4c07] <= 8'h14;
		memory[16'h4c08] <= 8'hfc;
		memory[16'h4c09] <= 8'h38;
		memory[16'h4c0a] <= 8'he3;
		memory[16'h4c0b] <= 8'h6e;
		memory[16'h4c0c] <= 8'h10;
		memory[16'h4c0d] <= 8'h66;
		memory[16'h4c0e] <= 8'h5c;
		memory[16'h4c0f] <= 8'h5e;
		memory[16'h4c10] <= 8'h26;
		memory[16'h4c11] <= 8'hd;
		memory[16'h4c12] <= 8'hcf;
		memory[16'h4c13] <= 8'h57;
		memory[16'h4c14] <= 8'hcd;
		memory[16'h4c15] <= 8'he6;
		memory[16'h4c16] <= 8'h94;
		memory[16'h4c17] <= 8'hfa;
		memory[16'h4c18] <= 8'h63;
		memory[16'h4c19] <= 8'h82;
		memory[16'h4c1a] <= 8'h7;
		memory[16'h4c1b] <= 8'h49;
		memory[16'h4c1c] <= 8'h93;
		memory[16'h4c1d] <= 8'ha6;
		memory[16'h4c1e] <= 8'hbb;
		memory[16'h4c1f] <= 8'he4;
		memory[16'h4c20] <= 8'h2f;
		memory[16'h4c21] <= 8'h68;
		memory[16'h4c22] <= 8'h8b;
		memory[16'h4c23] <= 8'h61;
		memory[16'h4c24] <= 8'h60;
		memory[16'h4c25] <= 8'hdf;
		memory[16'h4c26] <= 8'h76;
		memory[16'h4c27] <= 8'h5c;
		memory[16'h4c28] <= 8'h18;
		memory[16'h4c29] <= 8'h59;
		memory[16'h4c2a] <= 8'hca;
		memory[16'h4c2b] <= 8'h28;
		memory[16'h4c2c] <= 8'hc0;
		memory[16'h4c2d] <= 8'h27;
		memory[16'h4c2e] <= 8'h86;
		memory[16'h4c2f] <= 8'he6;
		memory[16'h4c30] <= 8'h34;
		memory[16'h4c31] <= 8'h55;
		memory[16'h4c32] <= 8'h3d;
		memory[16'h4c33] <= 8'h1;
		memory[16'h4c34] <= 8'h3c;
		memory[16'h4c35] <= 8'hd1;
		memory[16'h4c36] <= 8'hfb;
		memory[16'h4c37] <= 8'h9f;
		memory[16'h4c38] <= 8'h54;
		memory[16'h4c39] <= 8'h2;
		memory[16'h4c3a] <= 8'he8;
		memory[16'h4c3b] <= 8'he7;
		memory[16'h4c3c] <= 8'ha8;
		memory[16'h4c3d] <= 8'ha3;
		memory[16'h4c3e] <= 8'hcb;
		memory[16'h4c3f] <= 8'hd8;
		memory[16'h4c40] <= 8'hc;
		memory[16'h4c41] <= 8'h57;
		memory[16'h4c42] <= 8'h39;
		memory[16'h4c43] <= 8'h6c;
		memory[16'h4c44] <= 8'h36;
		memory[16'h4c45] <= 8'haf;
		memory[16'h4c46] <= 8'hc8;
		memory[16'h4c47] <= 8'h4e;
		memory[16'h4c48] <= 8'h9;
		memory[16'h4c49] <= 8'h92;
		memory[16'h4c4a] <= 8'h76;
		memory[16'h4c4b] <= 8'hc9;
		memory[16'h4c4c] <= 8'hb9;
		memory[16'h4c4d] <= 8'hfd;
		memory[16'h4c4e] <= 8'haf;
		memory[16'h4c4f] <= 8'hed;
		memory[16'h4c50] <= 8'h52;
		memory[16'h4c51] <= 8'hed;
		memory[16'h4c52] <= 8'hee;
		memory[16'h4c53] <= 8'h8e;
		memory[16'h4c54] <= 8'hbe;
		memory[16'h4c55] <= 8'he9;
		memory[16'h4c56] <= 8'h2d;
		memory[16'h4c57] <= 8'h12;
		memory[16'h4c58] <= 8'heb;
		memory[16'h4c59] <= 8'h15;
		memory[16'h4c5a] <= 8'hf9;
		memory[16'h4c5b] <= 8'h94;
		memory[16'h4c5c] <= 8'hb9;
		memory[16'h4c5d] <= 8'hc5;
		memory[16'h4c5e] <= 8'h6c;
		memory[16'h4c5f] <= 8'hc5;
		memory[16'h4c60] <= 8'h1c;
		memory[16'h4c61] <= 8'ha5;
		memory[16'h4c62] <= 8'h31;
		memory[16'h4c63] <= 8'h52;
		memory[16'h4c64] <= 8'h55;
		memory[16'h4c65] <= 8'hf9;
		memory[16'h4c66] <= 8'ha1;
		memory[16'h4c67] <= 8'h5e;
		memory[16'h4c68] <= 8'h8b;
		memory[16'h4c69] <= 8'h17;
		memory[16'h4c6a] <= 8'h27;
		memory[16'h4c6b] <= 8'h45;
		memory[16'h4c6c] <= 8'h14;
		memory[16'h4c6d] <= 8'hd6;
		memory[16'h4c6e] <= 8'h32;
		memory[16'h4c6f] <= 8'h67;
		memory[16'h4c70] <= 8'hc3;
		memory[16'h4c71] <= 8'h21;
		memory[16'h4c72] <= 8'hf5;
		memory[16'h4c73] <= 8'h82;
		memory[16'h4c74] <= 8'ha;
		memory[16'h4c75] <= 8'h23;
		memory[16'h4c76] <= 8'h94;
		memory[16'h4c77] <= 8'hf6;
		memory[16'h4c78] <= 8'h38;
		memory[16'h4c79] <= 8'h8e;
		memory[16'h4c7a] <= 8'h8a;
		memory[16'h4c7b] <= 8'hf1;
		memory[16'h4c7c] <= 8'h53;
		memory[16'h4c7d] <= 8'hf6;
		memory[16'h4c7e] <= 8'hb6;
		memory[16'h4c7f] <= 8'h6f;
		memory[16'h4c80] <= 8'h9b;
		memory[16'h4c81] <= 8'he7;
		memory[16'h4c82] <= 8'hc1;
		memory[16'h4c83] <= 8'hf0;
		memory[16'h4c84] <= 8'he0;
		memory[16'h4c85] <= 8'h62;
		memory[16'h4c86] <= 8'h4e;
		memory[16'h4c87] <= 8'h6c;
		memory[16'h4c88] <= 8'h7a;
		memory[16'h4c89] <= 8'h75;
		memory[16'h4c8a] <= 8'hb1;
		memory[16'h4c8b] <= 8'h8e;
		memory[16'h4c8c] <= 8'h4c;
		memory[16'h4c8d] <= 8'he3;
		memory[16'h4c8e] <= 8'hf5;
		memory[16'h4c8f] <= 8'hf;
		memory[16'h4c90] <= 8'h4;
		memory[16'h4c91] <= 8'heb;
		memory[16'h4c92] <= 8'h91;
		memory[16'h4c93] <= 8'hf;
		memory[16'h4c94] <= 8'he;
		memory[16'h4c95] <= 8'h26;
		memory[16'h4c96] <= 8'h5;
		memory[16'h4c97] <= 8'h46;
		memory[16'h4c98] <= 8'hb4;
		memory[16'h4c99] <= 8'h8f;
		memory[16'h4c9a] <= 8'h38;
		memory[16'h4c9b] <= 8'h7;
		memory[16'h4c9c] <= 8'h85;
		memory[16'h4c9d] <= 8'hee;
		memory[16'h4c9e] <= 8'h76;
		memory[16'h4c9f] <= 8'h20;
		memory[16'h4ca0] <= 8'hd6;
		memory[16'h4ca1] <= 8'h37;
		memory[16'h4ca2] <= 8'h11;
		memory[16'h4ca3] <= 8'hb6;
		memory[16'h4ca4] <= 8'h9a;
		memory[16'h4ca5] <= 8'h5f;
		memory[16'h4ca6] <= 8'h22;
		memory[16'h4ca7] <= 8'h14;
		memory[16'h4ca8] <= 8'hd5;
		memory[16'h4ca9] <= 8'hd3;
		memory[16'h4caa] <= 8'ha2;
		memory[16'h4cab] <= 8'h21;
		memory[16'h4cac] <= 8'hb7;
		memory[16'h4cad] <= 8'h98;
		memory[16'h4cae] <= 8'h30;
		memory[16'h4caf] <= 8'hbb;
		memory[16'h4cb0] <= 8'h83;
		memory[16'h4cb1] <= 8'hc2;
		memory[16'h4cb2] <= 8'hca;
		memory[16'h4cb3] <= 8'h91;
		memory[16'h4cb4] <= 8'he8;
		memory[16'h4cb5] <= 8'hcf;
		memory[16'h4cb6] <= 8'hd7;
		memory[16'h4cb7] <= 8'h9c;
		memory[16'h4cb8] <= 8'h5e;
		memory[16'h4cb9] <= 8'hf;
		memory[16'h4cba] <= 8'ha3;
		memory[16'h4cbb] <= 8'he3;
		memory[16'h4cbc] <= 8'hfe;
		memory[16'h4cbd] <= 8'h19;
		memory[16'h4cbe] <= 8'h4;
		memory[16'h4cbf] <= 8'hd4;
		memory[16'h4cc0] <= 8'h50;
		memory[16'h4cc1] <= 8'h15;
		memory[16'h4cc2] <= 8'h8a;
		memory[16'h4cc3] <= 8'hea;
		memory[16'h4cc4] <= 8'h74;
		memory[16'h4cc5] <= 8'had;
		memory[16'h4cc6] <= 8'hfe;
		memory[16'h4cc7] <= 8'h49;
		memory[16'h4cc8] <= 8'h80;
		memory[16'h4cc9] <= 8'ha1;
		memory[16'h4cca] <= 8'h6a;
		memory[16'h4ccb] <= 8'h37;
		memory[16'h4ccc] <= 8'h39;
		memory[16'h4ccd] <= 8'h9b;
		memory[16'h4cce] <= 8'hf3;
		memory[16'h4ccf] <= 8'hbc;
		memory[16'h4cd0] <= 8'h5d;
		memory[16'h4cd1] <= 8'hbd;
		memory[16'h4cd2] <= 8'h4d;
		memory[16'h4cd3] <= 8'h45;
		memory[16'h4cd4] <= 8'h8d;
		memory[16'h4cd5] <= 8'h24;
		memory[16'h4cd6] <= 8'he1;
		memory[16'h4cd7] <= 8'heb;
		memory[16'h4cd8] <= 8'h34;
		memory[16'h4cd9] <= 8'h84;
		memory[16'h4cda] <= 8'hcf;
		memory[16'h4cdb] <= 8'h32;
		memory[16'h4cdc] <= 8'h9d;
		memory[16'h4cdd] <= 8'hd3;
		memory[16'h4cde] <= 8'h6;
		memory[16'h4cdf] <= 8'hed;
		memory[16'h4ce0] <= 8'he8;
		memory[16'h4ce1] <= 8'h90;
		memory[16'h4ce2] <= 8'hd8;
		memory[16'h4ce3] <= 8'h5c;
		memory[16'h4ce4] <= 8'h3d;
		memory[16'h4ce5] <= 8'hd6;
		memory[16'h4ce6] <= 8'ha6;
		memory[16'h4ce7] <= 8'hbe;
		memory[16'h4ce8] <= 8'h77;
		memory[16'h4ce9] <= 8'h10;
		memory[16'h4cea] <= 8'hf5;
		memory[16'h4ceb] <= 8'hb0;
		memory[16'h4cec] <= 8'hab;
		memory[16'h4ced] <= 8'he8;
		memory[16'h4cee] <= 8'h6c;
		memory[16'h4cef] <= 8'h8;
		memory[16'h4cf0] <= 8'ha6;
		memory[16'h4cf1] <= 8'hb9;
		memory[16'h4cf2] <= 8'h4d;
		memory[16'h4cf3] <= 8'h33;
		memory[16'h4cf4] <= 8'hde;
		memory[16'h4cf5] <= 8'h2e;
		memory[16'h4cf6] <= 8'h1e;
		memory[16'h4cf7] <= 8'h12;
		memory[16'h4cf8] <= 8'hb2;
		memory[16'h4cf9] <= 8'hed;
		memory[16'h4cfa] <= 8'h44;
		memory[16'h4cfb] <= 8'h4f;
		memory[16'h4cfc] <= 8'hc0;
		memory[16'h4cfd] <= 8'h4a;
		memory[16'h4cfe] <= 8'h3d;
		memory[16'h4cff] <= 8'ha8;
		memory[16'h4d00] <= 8'hda;
		memory[16'h4d01] <= 8'h15;
		memory[16'h4d02] <= 8'h5;
		memory[16'h4d03] <= 8'h18;
		memory[16'h4d04] <= 8'heb;
		memory[16'h4d05] <= 8'hab;
		memory[16'h4d06] <= 8'hd6;
		memory[16'h4d07] <= 8'h63;
		memory[16'h4d08] <= 8'hbb;
		memory[16'h4d09] <= 8'hcb;
		memory[16'h4d0a] <= 8'h13;
		memory[16'h4d0b] <= 8'h67;
		memory[16'h4d0c] <= 8'hb4;
		memory[16'h4d0d] <= 8'h80;
		memory[16'h4d0e] <= 8'h6f;
		memory[16'h4d0f] <= 8'h5a;
		memory[16'h4d10] <= 8'h39;
		memory[16'h4d11] <= 8'hbd;
		memory[16'h4d12] <= 8'h8d;
		memory[16'h4d13] <= 8'h17;
		memory[16'h4d14] <= 8'heb;
		memory[16'h4d15] <= 8'hab;
		memory[16'h4d16] <= 8'h29;
		memory[16'h4d17] <= 8'h9e;
		memory[16'h4d18] <= 8'h99;
		memory[16'h4d19] <= 8'h6d;
		memory[16'h4d1a] <= 8'hed;
		memory[16'h4d1b] <= 8'h59;
		memory[16'h4d1c] <= 8'hb7;
		memory[16'h4d1d] <= 8'h2a;
		memory[16'h4d1e] <= 8'h2;
		memory[16'h4d1f] <= 8'h92;
		memory[16'h4d20] <= 8'h3f;
		memory[16'h4d21] <= 8'h7;
		memory[16'h4d22] <= 8'haa;
		memory[16'h4d23] <= 8'h2b;
		memory[16'h4d24] <= 8'hb2;
		memory[16'h4d25] <= 8'h80;
		memory[16'h4d26] <= 8'h8e;
		memory[16'h4d27] <= 8'h6d;
		memory[16'h4d28] <= 8'h4b;
		memory[16'h4d29] <= 8'ha1;
		memory[16'h4d2a] <= 8'hd4;
		memory[16'h4d2b] <= 8'hff;
		memory[16'h4d2c] <= 8'h21;
		memory[16'h4d2d] <= 8'h44;
		memory[16'h4d2e] <= 8'h59;
		memory[16'h4d2f] <= 8'h5b;
		memory[16'h4d30] <= 8'h1;
		memory[16'h4d31] <= 8'he6;
		memory[16'h4d32] <= 8'h72;
		memory[16'h4d33] <= 8'hec;
		memory[16'h4d34] <= 8'h92;
		memory[16'h4d35] <= 8'h9c;
		memory[16'h4d36] <= 8'h8a;
		memory[16'h4d37] <= 8'h2b;
		memory[16'h4d38] <= 8'h9;
		memory[16'h4d39] <= 8'h78;
		memory[16'h4d3a] <= 8'h84;
		memory[16'h4d3b] <= 8'hc1;
		memory[16'h4d3c] <= 8'ha2;
		memory[16'h4d3d] <= 8'h86;
		memory[16'h4d3e] <= 8'h53;
		memory[16'h4d3f] <= 8'he2;
		memory[16'h4d40] <= 8'h8d;
		memory[16'h4d41] <= 8'hfd;
		memory[16'h4d42] <= 8'hd;
		memory[16'h4d43] <= 8'h3f;
		memory[16'h4d44] <= 8'h7d;
		memory[16'h4d45] <= 8'h9b;
		memory[16'h4d46] <= 8'had;
		memory[16'h4d47] <= 8'hc8;
		memory[16'h4d48] <= 8'h3c;
		memory[16'h4d49] <= 8'h81;
		memory[16'h4d4a] <= 8'hc8;
		memory[16'h4d4b] <= 8'h5e;
		memory[16'h4d4c] <= 8'hc5;
		memory[16'h4d4d] <= 8'h21;
		memory[16'h4d4e] <= 8'hb9;
		memory[16'h4d4f] <= 8'hc6;
		memory[16'h4d50] <= 8'h8;
		memory[16'h4d51] <= 8'h2b;
		memory[16'h4d52] <= 8'hb3;
		memory[16'h4d53] <= 8'h9a;
		memory[16'h4d54] <= 8'hc7;
		memory[16'h4d55] <= 8'h3d;
		memory[16'h4d56] <= 8'hc5;
		memory[16'h4d57] <= 8'hd1;
		memory[16'h4d58] <= 8'hb5;
		memory[16'h4d59] <= 8'h49;
		memory[16'h4d5a] <= 8'h92;
		memory[16'h4d5b] <= 8'h58;
		memory[16'h4d5c] <= 8'hd0;
		memory[16'h4d5d] <= 8'he5;
		memory[16'h4d5e] <= 8'h3a;
		memory[16'h4d5f] <= 8'h5d;
		memory[16'h4d60] <= 8'he2;
		memory[16'h4d61] <= 8'h47;
		memory[16'h4d62] <= 8'h9d;
		memory[16'h4d63] <= 8'h5f;
		memory[16'h4d64] <= 8'he2;
		memory[16'h4d65] <= 8'h4a;
		memory[16'h4d66] <= 8'h27;
		memory[16'h4d67] <= 8'h1e;
		memory[16'h4d68] <= 8'hcb;
		memory[16'h4d69] <= 8'hef;
		memory[16'h4d6a] <= 8'h7c;
		memory[16'h4d6b] <= 8'h91;
		memory[16'h4d6c] <= 8'h11;
		memory[16'h4d6d] <= 8'h35;
		memory[16'h4d6e] <= 8'h57;
		memory[16'h4d6f] <= 8'h19;
		memory[16'h4d70] <= 8'h61;
		memory[16'h4d71] <= 8'ha;
		memory[16'h4d72] <= 8'hb3;
		memory[16'h4d73] <= 8'h28;
		memory[16'h4d74] <= 8'h48;
		memory[16'h4d75] <= 8'h78;
		memory[16'h4d76] <= 8'hf9;
		memory[16'h4d77] <= 8'hfd;
		memory[16'h4d78] <= 8'hc1;
		memory[16'h4d79] <= 8'h8b;
		memory[16'h4d7a] <= 8'h55;
		memory[16'h4d7b] <= 8'h91;
		memory[16'h4d7c] <= 8'h70;
		memory[16'h4d7d] <= 8'h8f;
		memory[16'h4d7e] <= 8'hef;
		memory[16'h4d7f] <= 8'h52;
		memory[16'h4d80] <= 8'hd6;
		memory[16'h4d81] <= 8'h8c;
		memory[16'h4d82] <= 8'hb1;
		memory[16'h4d83] <= 8'hb8;
		memory[16'h4d84] <= 8'hd6;
		memory[16'h4d85] <= 8'hd9;
		memory[16'h4d86] <= 8'hd7;
		memory[16'h4d87] <= 8'ha1;
		memory[16'h4d88] <= 8'hc8;
		memory[16'h4d89] <= 8'h53;
		memory[16'h4d8a] <= 8'h32;
		memory[16'h4d8b] <= 8'hd9;
		memory[16'h4d8c] <= 8'h89;
		memory[16'h4d8d] <= 8'h8a;
		memory[16'h4d8e] <= 8'hf2;
		memory[16'h4d8f] <= 8'hea;
		memory[16'h4d90] <= 8'h94;
		memory[16'h4d91] <= 8'ha5;
		memory[16'h4d92] <= 8'h12;
		memory[16'h4d93] <= 8'hdc;
		memory[16'h4d94] <= 8'h1d;
		memory[16'h4d95] <= 8'hc;
		memory[16'h4d96] <= 8'hda;
		memory[16'h4d97] <= 8'hdf;
		memory[16'h4d98] <= 8'h97;
		memory[16'h4d99] <= 8'h2f;
		memory[16'h4d9a] <= 8'h70;
		memory[16'h4d9b] <= 8'h8;
		memory[16'h4d9c] <= 8'hbf;
		memory[16'h4d9d] <= 8'h5f;
		memory[16'h4d9e] <= 8'h5a;
		memory[16'h4d9f] <= 8'h95;
		memory[16'h4da0] <= 8'heb;
		memory[16'h4da1] <= 8'hc;
		memory[16'h4da2] <= 8'h4e;
		memory[16'h4da3] <= 8'hc1;
		memory[16'h4da4] <= 8'he5;
		memory[16'h4da5] <= 8'h25;
		memory[16'h4da6] <= 8'h63;
		memory[16'h4da7] <= 8'had;
		memory[16'h4da8] <= 8'h78;
		memory[16'h4da9] <= 8'h95;
		memory[16'h4daa] <= 8'h87;
		memory[16'h4dab] <= 8'h1;
		memory[16'h4dac] <= 8'h1f;
		memory[16'h4dad] <= 8'h79;
		memory[16'h4dae] <= 8'heb;
		memory[16'h4daf] <= 8'hb4;
		memory[16'h4db0] <= 8'h1f;
		memory[16'h4db1] <= 8'hfe;
		memory[16'h4db2] <= 8'h90;
		memory[16'h4db3] <= 8'h3c;
		memory[16'h4db4] <= 8'ha;
		memory[16'h4db5] <= 8'h6a;
		memory[16'h4db6] <= 8'h1b;
		memory[16'h4db7] <= 8'ha1;
		memory[16'h4db8] <= 8'h9a;
		memory[16'h4db9] <= 8'h8c;
		memory[16'h4dba] <= 8'ha9;
		memory[16'h4dbb] <= 8'h59;
		memory[16'h4dbc] <= 8'heb;
		memory[16'h4dbd] <= 8'h4;
		memory[16'h4dbe] <= 8'hee;
		memory[16'h4dbf] <= 8'hd7;
		memory[16'h4dc0] <= 8'h10;
		memory[16'h4dc1] <= 8'h3c;
		memory[16'h4dc2] <= 8'h98;
		memory[16'h4dc3] <= 8'hf5;
		memory[16'h4dc4] <= 8'h61;
		memory[16'h4dc5] <= 8'hfb;
		memory[16'h4dc6] <= 8'ha2;
		memory[16'h4dc7] <= 8'hda;
		memory[16'h4dc8] <= 8'h91;
		memory[16'h4dc9] <= 8'h29;
		memory[16'h4dca] <= 8'hdb;
		memory[16'h4dcb] <= 8'hb0;
		memory[16'h4dcc] <= 8'ha3;
		memory[16'h4dcd] <= 8'hc7;
		memory[16'h4dce] <= 8'h64;
		memory[16'h4dcf] <= 8'hc2;
		memory[16'h4dd0] <= 8'hc5;
		memory[16'h4dd1] <= 8'hf5;
		memory[16'h4dd2] <= 8'hfe;
		memory[16'h4dd3] <= 8'hcf;
		memory[16'h4dd4] <= 8'h5f;
		memory[16'h4dd5] <= 8'h1a;
		memory[16'h4dd6] <= 8'h70;
		memory[16'h4dd7] <= 8'hf9;
		memory[16'h4dd8] <= 8'ha6;
		memory[16'h4dd9] <= 8'h1a;
		memory[16'h4dda] <= 8'h52;
		memory[16'h4ddb] <= 8'h91;
		memory[16'h4ddc] <= 8'h1e;
		memory[16'h4ddd] <= 8'h41;
		memory[16'h4dde] <= 8'h68;
		memory[16'h4ddf] <= 8'h2e;
		memory[16'h4de0] <= 8'h7d;
		memory[16'h4de1] <= 8'h1;
		memory[16'h4de2] <= 8'h23;
		memory[16'h4de3] <= 8'hdf;
		memory[16'h4de4] <= 8'hfc;
		memory[16'h4de5] <= 8'hc5;
		memory[16'h4de6] <= 8'hb9;
		memory[16'h4de7] <= 8'h8d;
		memory[16'h4de8] <= 8'hef;
		memory[16'h4de9] <= 8'h94;
		memory[16'h4dea] <= 8'h3e;
		memory[16'h4deb] <= 8'h92;
		memory[16'h4dec] <= 8'h5b;
		memory[16'h4ded] <= 8'ha2;
		memory[16'h4dee] <= 8'h54;
		memory[16'h4def] <= 8'h20;
		memory[16'h4df0] <= 8'h97;
		memory[16'h4df1] <= 8'h52;
		memory[16'h4df2] <= 8'hef;
		memory[16'h4df3] <= 8'hf7;
		memory[16'h4df4] <= 8'h6c;
		memory[16'h4df5] <= 8'h60;
		memory[16'h4df6] <= 8'hf0;
		memory[16'h4df7] <= 8'h12;
		memory[16'h4df8] <= 8'h7a;
		memory[16'h4df9] <= 8'h43;
		memory[16'h4dfa] <= 8'ha4;
		memory[16'h4dfb] <= 8'h98;
		memory[16'h4dfc] <= 8'h84;
		memory[16'h4dfd] <= 8'hc;
		memory[16'h4dfe] <= 8'hc6;
		memory[16'h4dff] <= 8'h1;
		memory[16'h4e00] <= 8'hd;
		memory[16'h4e01] <= 8'he9;
		memory[16'h4e02] <= 8'he0;
		memory[16'h4e03] <= 8'ha;
		memory[16'h4e04] <= 8'hae;
		memory[16'h4e05] <= 8'h99;
		memory[16'h4e06] <= 8'h97;
		memory[16'h4e07] <= 8'h9d;
		memory[16'h4e08] <= 8'h2e;
		memory[16'h4e09] <= 8'hd5;
		memory[16'h4e0a] <= 8'h2f;
		memory[16'h4e0b] <= 8'h89;
		memory[16'h4e0c] <= 8'h78;
		memory[16'h4e0d] <= 8'h83;
		memory[16'h4e0e] <= 8'haa;
		memory[16'h4e0f] <= 8'hf;
		memory[16'h4e10] <= 8'hd6;
		memory[16'h4e11] <= 8'h99;
		memory[16'h4e12] <= 8'h6;
		memory[16'h4e13] <= 8'h42;
		memory[16'h4e14] <= 8'hf9;
		memory[16'h4e15] <= 8'hf7;
		memory[16'h4e16] <= 8'h55;
		memory[16'h4e17] <= 8'h73;
		memory[16'h4e18] <= 8'h3a;
		memory[16'h4e19] <= 8'hf9;
		memory[16'h4e1a] <= 8'hb;
		memory[16'h4e1b] <= 8'hbe;
		memory[16'h4e1c] <= 8'h5;
		memory[16'h4e1d] <= 8'hd1;
		memory[16'h4e1e] <= 8'hbf;
		memory[16'h4e1f] <= 8'h13;
		memory[16'h4e20] <= 8'hba;
		memory[16'h4e21] <= 8'ha0;
		memory[16'h4e22] <= 8'h1d;
		memory[16'h4e23] <= 8'h69;
		memory[16'h4e24] <= 8'h39;
		memory[16'h4e25] <= 8'hb4;
		memory[16'h4e26] <= 8'h6;
		memory[16'h4e27] <= 8'h67;
		memory[16'h4e28] <= 8'h8a;
		memory[16'h4e29] <= 8'h36;
		memory[16'h4e2a] <= 8'hf1;
		memory[16'h4e2b] <= 8'h2;
		memory[16'h4e2c] <= 8'hb9;
		memory[16'h4e2d] <= 8'h9b;
		memory[16'h4e2e] <= 8'h11;
		memory[16'h4e2f] <= 8'h8f;
		memory[16'h4e30] <= 8'h34;
		memory[16'h4e31] <= 8'h18;
		memory[16'h4e32] <= 8'hd2;
		memory[16'h4e33] <= 8'h2e;
		memory[16'h4e34] <= 8'hf;
		memory[16'h4e35] <= 8'h27;
		memory[16'h4e36] <= 8'ha1;
		memory[16'h4e37] <= 8'h49;
		memory[16'h4e38] <= 8'h20;
		memory[16'h4e39] <= 8'had;
		memory[16'h4e3a] <= 8'h7;
		memory[16'h4e3b] <= 8'h25;
		memory[16'h4e3c] <= 8'h7e;
		memory[16'h4e3d] <= 8'hc6;
		memory[16'h4e3e] <= 8'h38;
		memory[16'h4e3f] <= 8'h39;
		memory[16'h4e40] <= 8'h66;
		memory[16'h4e41] <= 8'h55;
		memory[16'h4e42] <= 8'ha2;
		memory[16'h4e43] <= 8'ha0;
		memory[16'h4e44] <= 8'ha;
		memory[16'h4e45] <= 8'ha8;
		memory[16'h4e46] <= 8'h7;
		memory[16'h4e47] <= 8'h94;
		memory[16'h4e48] <= 8'hde;
		memory[16'h4e49] <= 8'hf8;
		memory[16'h4e4a] <= 8'h96;
		memory[16'h4e4b] <= 8'h98;
		memory[16'h4e4c] <= 8'h93;
		memory[16'h4e4d] <= 8'ha7;
		memory[16'h4e4e] <= 8'h27;
		memory[16'h4e4f] <= 8'hc8;
		memory[16'h4e50] <= 8'hbf;
		memory[16'h4e51] <= 8'hf9;
		memory[16'h4e52] <= 8'hf6;
		memory[16'h4e53] <= 8'hce;
		memory[16'h4e54] <= 8'h20;
		memory[16'h4e55] <= 8'h97;
		memory[16'h4e56] <= 8'h17;
		memory[16'h4e57] <= 8'h40;
		memory[16'h4e58] <= 8'h44;
		memory[16'h4e59] <= 8'h1e;
		memory[16'h4e5a] <= 8'h66;
		memory[16'h4e5b] <= 8'hc3;
		memory[16'h4e5c] <= 8'he5;
		memory[16'h4e5d] <= 8'h9e;
		memory[16'h4e5e] <= 8'hfc;
		memory[16'h4e5f] <= 8'h4b;
		memory[16'h4e60] <= 8'hf4;
		memory[16'h4e61] <= 8'h9e;
		memory[16'h4e62] <= 8'heb;
		memory[16'h4e63] <= 8'hfe;
		memory[16'h4e64] <= 8'h46;
		memory[16'h4e65] <= 8'hf3;
		memory[16'h4e66] <= 8'h92;
		memory[16'h4e67] <= 8'h25;
		memory[16'h4e68] <= 8'heb;
		memory[16'h4e69] <= 8'h28;
		memory[16'h4e6a] <= 8'hbd;
		memory[16'h4e6b] <= 8'h7f;
		memory[16'h4e6c] <= 8'hcf;
		memory[16'h4e6d] <= 8'he4;
		memory[16'h4e6e] <= 8'h47;
		memory[16'h4e6f] <= 8'h8f;
		memory[16'h4e70] <= 8'hde;
		memory[16'h4e71] <= 8'h3d;
		memory[16'h4e72] <= 8'h5d;
		memory[16'h4e73] <= 8'hfe;
		memory[16'h4e74] <= 8'hd4;
		memory[16'h4e75] <= 8'h75;
		memory[16'h4e76] <= 8'h3f;
		memory[16'h4e77] <= 8'h19;
		memory[16'h4e78] <= 8'h93;
		memory[16'h4e79] <= 8'ha5;
		memory[16'h4e7a] <= 8'hdc;
		memory[16'h4e7b] <= 8'h78;
		memory[16'h4e7c] <= 8'h43;
		memory[16'h4e7d] <= 8'hd8;
		memory[16'h4e7e] <= 8'hc4;
		memory[16'h4e7f] <= 8'h37;
		memory[16'h4e80] <= 8'h76;
		memory[16'h4e81] <= 8'haf;
		memory[16'h4e82] <= 8'h35;
		memory[16'h4e83] <= 8'hbc;
		memory[16'h4e84] <= 8'ha2;
		memory[16'h4e85] <= 8'hc7;
		memory[16'h4e86] <= 8'he1;
		memory[16'h4e87] <= 8'h8e;
		memory[16'h4e88] <= 8'hef;
		memory[16'h4e89] <= 8'h9e;
		memory[16'h4e8a] <= 8'hd;
		memory[16'h4e8b] <= 8'hbf;
		memory[16'h4e8c] <= 8'h83;
		memory[16'h4e8d] <= 8'h54;
		memory[16'h4e8e] <= 8'h4e;
		memory[16'h4e8f] <= 8'h61;
		memory[16'h4e90] <= 8'h91;
		memory[16'h4e91] <= 8'hab;
		memory[16'h4e92] <= 8'h5f;
		memory[16'h4e93] <= 8'h65;
		memory[16'h4e94] <= 8'h20;
		memory[16'h4e95] <= 8'h9e;
		memory[16'h4e96] <= 8'h7e;
		memory[16'h4e97] <= 8'hb4;
		memory[16'h4e98] <= 8'h43;
		memory[16'h4e99] <= 8'h5a;
		memory[16'h4e9a] <= 8'h2c;
		memory[16'h4e9b] <= 8'h87;
		memory[16'h4e9c] <= 8'h32;
		memory[16'h4e9d] <= 8'hf0;
		memory[16'h4e9e] <= 8'hbe;
		memory[16'h4e9f] <= 8'ha8;
		memory[16'h4ea0] <= 8'ha0;
		memory[16'h4ea1] <= 8'hf4;
		memory[16'h4ea2] <= 8'h65;
		memory[16'h4ea3] <= 8'h42;
		memory[16'h4ea4] <= 8'hbb;
		memory[16'h4ea5] <= 8'h46;
		memory[16'h4ea6] <= 8'hd0;
		memory[16'h4ea7] <= 8'hab;
		memory[16'h4ea8] <= 8'he5;
		memory[16'h4ea9] <= 8'hdd;
		memory[16'h4eaa] <= 8'h6a;
		memory[16'h4eab] <= 8'h68;
		memory[16'h4eac] <= 8'h31;
		memory[16'h4ead] <= 8'hb8;
		memory[16'h4eae] <= 8'hc9;
		memory[16'h4eaf] <= 8'hc2;
		memory[16'h4eb0] <= 8'h63;
		memory[16'h4eb1] <= 8'h28;
		memory[16'h4eb2] <= 8'h28;
		memory[16'h4eb3] <= 8'h84;
		memory[16'h4eb4] <= 8'hc7;
		memory[16'h4eb5] <= 8'ha6;
		memory[16'h4eb6] <= 8'h38;
		memory[16'h4eb7] <= 8'ha;
		memory[16'h4eb8] <= 8'h1;
		memory[16'h4eb9] <= 8'h64;
		memory[16'h4eba] <= 8'h91;
		memory[16'h4ebb] <= 8'h33;
		memory[16'h4ebc] <= 8'h55;
		memory[16'h4ebd] <= 8'h50;
		memory[16'h4ebe] <= 8'hdc;
		memory[16'h4ebf] <= 8'hf5;
		memory[16'h4ec0] <= 8'h44;
		memory[16'h4ec1] <= 8'h41;
		memory[16'h4ec2] <= 8'h37;
		memory[16'h4ec3] <= 8'hff;
		memory[16'h4ec4] <= 8'h87;
		memory[16'h4ec5] <= 8'h8;
		memory[16'h4ec6] <= 8'haa;
		memory[16'h4ec7] <= 8'h6c;
		memory[16'h4ec8] <= 8'he5;
		memory[16'h4ec9] <= 8'h14;
		memory[16'h4eca] <= 8'hd4;
		memory[16'h4ecb] <= 8'h17;
		memory[16'h4ecc] <= 8'hcc;
		memory[16'h4ecd] <= 8'h9d;
		memory[16'h4ece] <= 8'hd9;
		memory[16'h4ecf] <= 8'h30;
		memory[16'h4ed0] <= 8'hc6;
		memory[16'h4ed1] <= 8'h1;
		memory[16'h4ed2] <= 8'hb4;
		memory[16'h4ed3] <= 8'h8d;
		memory[16'h4ed4] <= 8'ha8;
		memory[16'h4ed5] <= 8'hec;
		memory[16'h4ed6] <= 8'h97;
		memory[16'h4ed7] <= 8'ha9;
		memory[16'h4ed8] <= 8'h50;
		memory[16'h4ed9] <= 8'h29;
		memory[16'h4eda] <= 8'hdc;
		memory[16'h4edb] <= 8'ha5;
		memory[16'h4edc] <= 8'h79;
		memory[16'h4edd] <= 8'hb8;
		memory[16'h4ede] <= 8'h9a;
		memory[16'h4edf] <= 8'hbd;
		memory[16'h4ee0] <= 8'hf9;
		memory[16'h4ee1] <= 8'hd2;
		memory[16'h4ee2] <= 8'hbc;
		memory[16'h4ee3] <= 8'h81;
		memory[16'h4ee4] <= 8'hda;
		memory[16'h4ee5] <= 8'h67;
		memory[16'h4ee6] <= 8'hed;
		memory[16'h4ee7] <= 8'hbf;
		memory[16'h4ee8] <= 8'h7b;
		memory[16'h4ee9] <= 8'hc2;
		memory[16'h4eea] <= 8'hd6;
		memory[16'h4eeb] <= 8'h48;
		memory[16'h4eec] <= 8'h5f;
		memory[16'h4eed] <= 8'hb0;
		memory[16'h4eee] <= 8'h78;
		memory[16'h4eef] <= 8'h25;
		memory[16'h4ef0] <= 8'hb1;
		memory[16'h4ef1] <= 8'h2c;
		memory[16'h4ef2] <= 8'hb2;
		memory[16'h4ef3] <= 8'h59;
		memory[16'h4ef4] <= 8'h18;
		memory[16'h4ef5] <= 8'h4a;
		memory[16'h4ef6] <= 8'h2;
		memory[16'h4ef7] <= 8'h68;
		memory[16'h4ef8] <= 8'h73;
		memory[16'h4ef9] <= 8'hdf;
		memory[16'h4efa] <= 8'he;
		memory[16'h4efb] <= 8'hec;
		memory[16'h4efc] <= 8'h97;
		memory[16'h4efd] <= 8'ha8;
		memory[16'h4efe] <= 8'ha9;
		memory[16'h4eff] <= 8'h91;
		memory[16'h4f00] <= 8'h7a;
		memory[16'h4f01] <= 8'h65;
		memory[16'h4f02] <= 8'h12;
		memory[16'h4f03] <= 8'h54;
		memory[16'h4f04] <= 8'hcc;
		memory[16'h4f05] <= 8'hff;
		memory[16'h4f06] <= 8'h14;
		memory[16'h4f07] <= 8'h48;
		memory[16'h4f08] <= 8'hc1;
		memory[16'h4f09] <= 8'hea;
		memory[16'h4f0a] <= 8'h90;
		memory[16'h4f0b] <= 8'h21;
		memory[16'h4f0c] <= 8'h9a;
		memory[16'h4f0d] <= 8'h8;
		memory[16'h4f0e] <= 8'h46;
		memory[16'h4f0f] <= 8'h4c;
		memory[16'h4f10] <= 8'h34;
		memory[16'h4f11] <= 8'hf9;
		memory[16'h4f12] <= 8'ha5;
		memory[16'h4f13] <= 8'h4c;
		memory[16'h4f14] <= 8'h43;
		memory[16'h4f15] <= 8'ha8;
		memory[16'h4f16] <= 8'hb4;
		memory[16'h4f17] <= 8'hb6;
		memory[16'h4f18] <= 8'h87;
		memory[16'h4f19] <= 8'hc2;
		memory[16'h4f1a] <= 8'ha2;
		memory[16'h4f1b] <= 8'h1e;
		memory[16'h4f1c] <= 8'h6b;
		memory[16'h4f1d] <= 8'h4b;
		memory[16'h4f1e] <= 8'haf;
		memory[16'h4f1f] <= 8'he5;
		memory[16'h4f20] <= 8'hb0;
		memory[16'h4f21] <= 8'hc1;
		memory[16'h4f22] <= 8'h3a;
		memory[16'h4f23] <= 8'h7d;
		memory[16'h4f24] <= 8'hc1;
		memory[16'h4f25] <= 8'h4e;
		memory[16'h4f26] <= 8'hc5;
		memory[16'h4f27] <= 8'h82;
		memory[16'h4f28] <= 8'h38;
		memory[16'h4f29] <= 8'h55;
		memory[16'h4f2a] <= 8'ha3;
		memory[16'h4f2b] <= 8'hd3;
		memory[16'h4f2c] <= 8'h5d;
		memory[16'h4f2d] <= 8'hea;
		memory[16'h4f2e] <= 8'h1f;
		memory[16'h4f2f] <= 8'h91;
		memory[16'h4f30] <= 8'he3;
		memory[16'h4f31] <= 8'hc4;
		memory[16'h4f32] <= 8'hdd;
		memory[16'h4f33] <= 8'h26;
		memory[16'h4f34] <= 8'h6c;
		memory[16'h4f35] <= 8'h91;
		memory[16'h4f36] <= 8'hdc;
		memory[16'h4f37] <= 8'hf3;
		memory[16'h4f38] <= 8'h54;
		memory[16'h4f39] <= 8'h7e;
		memory[16'h4f3a] <= 8'h12;
		memory[16'h4f3b] <= 8'hbf;
		memory[16'h4f3c] <= 8'hc9;
		memory[16'h4f3d] <= 8'hc1;
		memory[16'h4f3e] <= 8'ha4;
		memory[16'h4f3f] <= 8'h79;
		memory[16'h4f40] <= 8'h83;
		memory[16'h4f41] <= 8'hde;
		memory[16'h4f42] <= 8'hf6;
		memory[16'h4f43] <= 8'h44;
		memory[16'h4f44] <= 8'h2c;
		memory[16'h4f45] <= 8'hbb;
		memory[16'h4f46] <= 8'hc6;
		memory[16'h4f47] <= 8'h65;
		memory[16'h4f48] <= 8'h10;
		memory[16'h4f49] <= 8'h6a;
		memory[16'h4f4a] <= 8'h38;
		memory[16'h4f4b] <= 8'h6d;
		memory[16'h4f4c] <= 8'h54;
		memory[16'h4f4d] <= 8'h57;
		memory[16'h4f4e] <= 8'hfe;
		memory[16'h4f4f] <= 8'h37;
		memory[16'h4f50] <= 8'h1b;
		memory[16'h4f51] <= 8'hdb;
		memory[16'h4f52] <= 8'h5d;
		memory[16'h4f53] <= 8'h88;
		memory[16'h4f54] <= 8'h6d;
		memory[16'h4f55] <= 8'h39;
		memory[16'h4f56] <= 8'h7b;
		memory[16'h4f57] <= 8'hc1;
		memory[16'h4f58] <= 8'hb7;
		memory[16'h4f59] <= 8'h8d;
		memory[16'h4f5a] <= 8'h80;
		memory[16'h4f5b] <= 8'h80;
		memory[16'h4f5c] <= 8'h4f;
		memory[16'h4f5d] <= 8'h24;
		memory[16'h4f5e] <= 8'hf9;
		memory[16'h4f5f] <= 8'hd2;
		memory[16'h4f60] <= 8'h3;
		memory[16'h4f61] <= 8'hf0;
		memory[16'h4f62] <= 8'h16;
		memory[16'h4f63] <= 8'h2f;
		memory[16'h4f64] <= 8'hab;
		memory[16'h4f65] <= 8'hdc;
		memory[16'h4f66] <= 8'h94;
		memory[16'h4f67] <= 8'hbc;
		memory[16'h4f68] <= 8'h46;
		memory[16'h4f69] <= 8'hcc;
		memory[16'h4f6a] <= 8'h29;
		memory[16'h4f6b] <= 8'h9a;
		memory[16'h4f6c] <= 8'h23;
		memory[16'h4f6d] <= 8'h28;
		memory[16'h4f6e] <= 8'hd1;
		memory[16'h4f6f] <= 8'h3f;
		memory[16'h4f70] <= 8'h3;
		memory[16'h4f71] <= 8'h2e;
		memory[16'h4f72] <= 8'hc7;
		memory[16'h4f73] <= 8'h70;
		memory[16'h4f74] <= 8'h67;
		memory[16'h4f75] <= 8'h42;
		memory[16'h4f76] <= 8'h31;
		memory[16'h4f77] <= 8'h1e;
		memory[16'h4f78] <= 8'hd0;
		memory[16'h4f79] <= 8'hb1;
		memory[16'h4f7a] <= 8'h9e;
		memory[16'h4f7b] <= 8'h1f;
		memory[16'h4f7c] <= 8'hd6;
		memory[16'h4f7d] <= 8'h98;
		memory[16'h4f7e] <= 8'hf1;
		memory[16'h4f7f] <= 8'hd9;
		memory[16'h4f80] <= 8'h88;
		memory[16'h4f81] <= 8'h7;
		memory[16'h4f82] <= 8'h8;
		memory[16'h4f83] <= 8'h33;
		memory[16'h4f84] <= 8'he3;
		memory[16'h4f85] <= 8'h9d;
		memory[16'h4f86] <= 8'hef;
		memory[16'h4f87] <= 8'h2a;
		memory[16'h4f88] <= 8'h69;
		memory[16'h4f89] <= 8'h19;
		memory[16'h4f8a] <= 8'hc4;
		memory[16'h4f8b] <= 8'h8d;
		memory[16'h4f8c] <= 8'h41;
		memory[16'h4f8d] <= 8'h96;
		memory[16'h4f8e] <= 8'hcc;
		memory[16'h4f8f] <= 8'h44;
		memory[16'h4f90] <= 8'hc4;
		memory[16'h4f91] <= 8'h93;
		memory[16'h4f92] <= 8'hb5;
		memory[16'h4f93] <= 8'h2c;
		memory[16'h4f94] <= 8'hd5;
		memory[16'h4f95] <= 8'he6;
		memory[16'h4f96] <= 8'h4a;
		memory[16'h4f97] <= 8'ha5;
		memory[16'h4f98] <= 8'h98;
		memory[16'h4f99] <= 8'he9;
		memory[16'h4f9a] <= 8'hc4;
		memory[16'h4f9b] <= 8'h6e;
		memory[16'h4f9c] <= 8'h81;
		memory[16'h4f9d] <= 8'hb5;
		memory[16'h4f9e] <= 8'h47;
		memory[16'h4f9f] <= 8'h9;
		memory[16'h4fa0] <= 8'hbc;
		memory[16'h4fa1] <= 8'h4f;
		memory[16'h4fa2] <= 8'h3c;
		memory[16'h4fa3] <= 8'ha0;
		memory[16'h4fa4] <= 8'hec;
		memory[16'h4fa5] <= 8'h2c;
		memory[16'h4fa6] <= 8'hca;
		memory[16'h4fa7] <= 8'h56;
		memory[16'h4fa8] <= 8'h45;
		memory[16'h4fa9] <= 8'h8e;
		memory[16'h4faa] <= 8'he3;
		memory[16'h4fab] <= 8'h86;
		memory[16'h4fac] <= 8'h24;
		memory[16'h4fad] <= 8'haf;
		memory[16'h4fae] <= 8'hca;
		memory[16'h4faf] <= 8'he9;
		memory[16'h4fb0] <= 8'h42;
		memory[16'h4fb1] <= 8'h7f;
		memory[16'h4fb2] <= 8'h15;
		memory[16'h4fb3] <= 8'h17;
		memory[16'h4fb4] <= 8'h66;
		memory[16'h4fb5] <= 8'h5f;
		memory[16'h4fb6] <= 8'hbd;
		memory[16'h4fb7] <= 8'hfe;
		memory[16'h4fb8] <= 8'h48;
		memory[16'h4fb9] <= 8'h81;
		memory[16'h4fba] <= 8'h6c;
		memory[16'h4fbb] <= 8'hc9;
		memory[16'h4fbc] <= 8'h37;
		memory[16'h4fbd] <= 8'hb3;
		memory[16'h4fbe] <= 8'hd2;
		memory[16'h4fbf] <= 8'hf3;
		memory[16'h4fc0] <= 8'h2;
		memory[16'h4fc1] <= 8'hf;
		memory[16'h4fc2] <= 8'h93;
		memory[16'h4fc3] <= 8'hef;
		memory[16'h4fc4] <= 8'h3b;
		memory[16'h4fc5] <= 8'h5d;
		memory[16'h4fc6] <= 8'h45;
		memory[16'h4fc7] <= 8'h80;
		memory[16'h4fc8] <= 8'hec;
		memory[16'h4fc9] <= 8'h28;
		memory[16'h4fca] <= 8'h6;
		memory[16'h4fcb] <= 8'h10;
		memory[16'h4fcc] <= 8'hd7;
		memory[16'h4fcd] <= 8'hd0;
		memory[16'h4fce] <= 8'hf9;
		memory[16'h4fcf] <= 8'h19;
		memory[16'h4fd0] <= 8'h50;
		memory[16'h4fd1] <= 8'he;
		memory[16'h4fd2] <= 8'h30;
		memory[16'h4fd3] <= 8'hb6;
		memory[16'h4fd4] <= 8'h6e;
		memory[16'h4fd5] <= 8'hed;
		memory[16'h4fd6] <= 8'hb4;
		memory[16'h4fd7] <= 8'hb6;
		memory[16'h4fd8] <= 8'h6f;
		memory[16'h4fd9] <= 8'h20;
		memory[16'h4fda] <= 8'h80;
		memory[16'h4fdb] <= 8'ha6;
		memory[16'h4fdc] <= 8'hd3;
		memory[16'h4fdd] <= 8'h52;
		memory[16'h4fde] <= 8'h99;
		memory[16'h4fdf] <= 8'hd5;
		memory[16'h4fe0] <= 8'h61;
		memory[16'h4fe1] <= 8'h2d;
		memory[16'h4fe2] <= 8'hc4;
		memory[16'h4fe3] <= 8'h9c;
		memory[16'h4fe4] <= 8'h8a;
		memory[16'h4fe5] <= 8'h9;
		memory[16'h4fe6] <= 8'h1c;
		memory[16'h4fe7] <= 8'h76;
		memory[16'h4fe8] <= 8'h31;
		memory[16'h4fe9] <= 8'h22;
		memory[16'h4fea] <= 8'h87;
		memory[16'h4feb] <= 8'h8;
		memory[16'h4fec] <= 8'hf3;
		memory[16'h4fed] <= 8'h80;
		memory[16'h4fee] <= 8'h21;
		memory[16'h4fef] <= 8'h43;
		memory[16'h4ff0] <= 8'h8f;
		memory[16'h4ff1] <= 8'h52;
		memory[16'h4ff2] <= 8'hf9;
		memory[16'h4ff3] <= 8'hfd;
		memory[16'h4ff4] <= 8'h3f;
		memory[16'h4ff5] <= 8'had;
		memory[16'h4ff6] <= 8'hb3;
		memory[16'h4ff7] <= 8'hae;
		memory[16'h4ff8] <= 8'hcd;
		memory[16'h4ff9] <= 8'h33;
		memory[16'h4ffa] <= 8'h54;
		memory[16'h4ffb] <= 8'ha0;
		memory[16'h4ffc] <= 8'h86;
		memory[16'h4ffd] <= 8'hee;
		memory[16'h4ffe] <= 8'h75;
		memory[16'h4fff] <= 8'he7;
		memory[16'h5000] <= 8'h1b;
		memory[16'h5001] <= 8'h3a;
		memory[16'h5002] <= 8'h84;
		memory[16'h5003] <= 8'ha5;
		memory[16'h5004] <= 8'h43;
		memory[16'h5005] <= 8'ha0;
		memory[16'h5006] <= 8'h1c;
		memory[16'h5007] <= 8'h75;
		memory[16'h5008] <= 8'hc3;
		memory[16'h5009] <= 8'ha3;
		memory[16'h500a] <= 8'h7d;
		memory[16'h500b] <= 8'hb6;
		memory[16'h500c] <= 8'h23;
		memory[16'h500d] <= 8'h9f;
		memory[16'h500e] <= 8'hf9;
		memory[16'h500f] <= 8'hb2;
		memory[16'h5010] <= 8'hf1;
		memory[16'h5011] <= 8'hf2;
		memory[16'h5012] <= 8'haf;
		memory[16'h5013] <= 8'h30;
		memory[16'h5014] <= 8'h9f;
		memory[16'h5015] <= 8'h63;
		memory[16'h5016] <= 8'hdf;
		memory[16'h5017] <= 8'h6c;
		memory[16'h5018] <= 8'h96;
		memory[16'h5019] <= 8'h33;
		memory[16'h501a] <= 8'hc;
		memory[16'h501b] <= 8'h1c;
		memory[16'h501c] <= 8'h21;
		memory[16'h501d] <= 8'h81;
		memory[16'h501e] <= 8'h4;
		memory[16'h501f] <= 8'h3c;
		memory[16'h5020] <= 8'hbb;
		memory[16'h5021] <= 8'h88;
		memory[16'h5022] <= 8'he2;
		memory[16'h5023] <= 8'hff;
		memory[16'h5024] <= 8'h28;
		memory[16'h5025] <= 8'hfe;
		memory[16'h5026] <= 8'h74;
		memory[16'h5027] <= 8'heb;
		memory[16'h5028] <= 8'ha1;
		memory[16'h5029] <= 8'hf1;
		memory[16'h502a] <= 8'ha1;
		memory[16'h502b] <= 8'hc4;
		memory[16'h502c] <= 8'h90;
		memory[16'h502d] <= 8'h9a;
		memory[16'h502e] <= 8'h77;
		memory[16'h502f] <= 8'h81;
		memory[16'h5030] <= 8'h8c;
		memory[16'h5031] <= 8'h26;
		memory[16'h5032] <= 8'hb2;
		memory[16'h5033] <= 8'h2b;
		memory[16'h5034] <= 8'h89;
		memory[16'h5035] <= 8'h91;
		memory[16'h5036] <= 8'h97;
		memory[16'h5037] <= 8'h20;
		memory[16'h5038] <= 8'hc4;
		memory[16'h5039] <= 8'ha3;
		memory[16'h503a] <= 8'h3c;
		memory[16'h503b] <= 8'he6;
		memory[16'h503c] <= 8'h25;
		memory[16'h503d] <= 8'h40;
		memory[16'h503e] <= 8'h22;
		memory[16'h503f] <= 8'he0;
		memory[16'h5040] <= 8'hc8;
		memory[16'h5041] <= 8'h4;
		memory[16'h5042] <= 8'hdf;
		memory[16'h5043] <= 8'hf1;
		memory[16'h5044] <= 8'h2;
		memory[16'h5045] <= 8'h53;
		memory[16'h5046] <= 8'hdc;
		memory[16'h5047] <= 8'ha3;
		memory[16'h5048] <= 8'h45;
		memory[16'h5049] <= 8'h7e;
		memory[16'h504a] <= 8'h68;
		memory[16'h504b] <= 8'hd5;
		memory[16'h504c] <= 8'h18;
		memory[16'h504d] <= 8'hdf;
		memory[16'h504e] <= 8'h57;
		memory[16'h504f] <= 8'ha5;
		memory[16'h5050] <= 8'h5;
		memory[16'h5051] <= 8'h9;
		memory[16'h5052] <= 8'hd0;
		memory[16'h5053] <= 8'h8f;
		memory[16'h5054] <= 8'h9a;
		memory[16'h5055] <= 8'h68;
		memory[16'h5056] <= 8'haf;
		memory[16'h5057] <= 8'h5e;
		memory[16'h5058] <= 8'hb;
		memory[16'h5059] <= 8'heb;
		memory[16'h505a] <= 8'h44;
		memory[16'h505b] <= 8'h30;
		memory[16'h505c] <= 8'h2c;
		memory[16'h505d] <= 8'h67;
		memory[16'h505e] <= 8'h11;
		memory[16'h505f] <= 8'hf4;
		memory[16'h5060] <= 8'h6b;
		memory[16'h5061] <= 8'hf0;
		memory[16'h5062] <= 8'he5;
		memory[16'h5063] <= 8'h6e;
		memory[16'h5064] <= 8'h44;
		memory[16'h5065] <= 8'hc2;
		memory[16'h5066] <= 8'h11;
		memory[16'h5067] <= 8'h89;
		memory[16'h5068] <= 8'h40;
		memory[16'h5069] <= 8'h79;
		memory[16'h506a] <= 8'h5e;
		memory[16'h506b] <= 8'h58;
		memory[16'h506c] <= 8'h58;
		memory[16'h506d] <= 8'hb5;
		memory[16'h506e] <= 8'hfd;
		memory[16'h506f] <= 8'h5e;
		memory[16'h5070] <= 8'hbe;
		memory[16'h5071] <= 8'hce;
		memory[16'h5072] <= 8'hed;
		memory[16'h5073] <= 8'h58;
		memory[16'h5074] <= 8'h36;
		memory[16'h5075] <= 8'h9c;
		memory[16'h5076] <= 8'hb7;
		memory[16'h5077] <= 8'h41;
		memory[16'h5078] <= 8'h87;
		memory[16'h5079] <= 8'hfb;
		memory[16'h507a] <= 8'h72;
		memory[16'h507b] <= 8'hb3;
		memory[16'h507c] <= 8'h62;
		memory[16'h507d] <= 8'h83;
		memory[16'h507e] <= 8'ha8;
		memory[16'h507f] <= 8'hce;
		memory[16'h5080] <= 8'h73;
		memory[16'h5081] <= 8'h8d;
		memory[16'h5082] <= 8'h3c;
		memory[16'h5083] <= 8'hb7;
		memory[16'h5084] <= 8'h4f;
		memory[16'h5085] <= 8'h4d;
		memory[16'h5086] <= 8'h40;
		memory[16'h5087] <= 8'h8f;
		memory[16'h5088] <= 8'hc7;
		memory[16'h5089] <= 8'h9f;
		memory[16'h508a] <= 8'he8;
		memory[16'h508b] <= 8'h1f;
		memory[16'h508c] <= 8'h54;
		memory[16'h508d] <= 8'he5;
		memory[16'h508e] <= 8'h7d;
		memory[16'h508f] <= 8'h13;
		memory[16'h5090] <= 8'hb3;
		memory[16'h5091] <= 8'h6a;
		memory[16'h5092] <= 8'h6b;
		memory[16'h5093] <= 8'he9;
		memory[16'h5094] <= 8'h6;
		memory[16'h5095] <= 8'h22;
		memory[16'h5096] <= 8'h2b;
		memory[16'h5097] <= 8'h8e;
		memory[16'h5098] <= 8'h1e;
		memory[16'h5099] <= 8'h9d;
		memory[16'h509a] <= 8'h41;
		memory[16'h509b] <= 8'h80;
		memory[16'h509c] <= 8'h20;
		memory[16'h509d] <= 8'he9;
		memory[16'h509e] <= 8'h4e;
		memory[16'h509f] <= 8'h93;
		memory[16'h50a0] <= 8'h77;
		memory[16'h50a1] <= 8'h8a;
		memory[16'h50a2] <= 8'h4b;
		memory[16'h50a3] <= 8'hc6;
		memory[16'h50a4] <= 8'hd8;
		memory[16'h50a5] <= 8'h8b;
		memory[16'h50a6] <= 8'h56;
		memory[16'h50a7] <= 8'h9f;
		memory[16'h50a8] <= 8'h2a;
		memory[16'h50a9] <= 8'h3e;
		memory[16'h50aa] <= 8'hbe;
		memory[16'h50ab] <= 8'h7f;
		memory[16'h50ac] <= 8'h23;
		memory[16'h50ad] <= 8'h3c;
		memory[16'h50ae] <= 8'h92;
		memory[16'h50af] <= 8'hd7;
		memory[16'h50b0] <= 8'ha6;
		memory[16'h50b1] <= 8'hfd;
		memory[16'h50b2] <= 8'hc0;
		memory[16'h50b3] <= 8'had;
		memory[16'h50b4] <= 8'h20;
		memory[16'h50b5] <= 8'heb;
		memory[16'h50b6] <= 8'h3b;
		memory[16'h50b7] <= 8'h3e;
		memory[16'h50b8] <= 8'h88;
		memory[16'h50b9] <= 8'h7c;
		memory[16'h50ba] <= 8'hbe;
		memory[16'h50bb] <= 8'ha8;
		memory[16'h50bc] <= 8'h66;
		memory[16'h50bd] <= 8'hd;
		memory[16'h50be] <= 8'h3c;
		memory[16'h50bf] <= 8'hdd;
		memory[16'h50c0] <= 8'h97;
		memory[16'h50c1] <= 8'h87;
		memory[16'h50c2] <= 8'ha3;
		memory[16'h50c3] <= 8'h6f;
		memory[16'h50c4] <= 8'h12;
		memory[16'h50c5] <= 8'hf9;
		memory[16'h50c6] <= 8'he;
		memory[16'h50c7] <= 8'h3d;
		memory[16'h50c8] <= 8'h37;
		memory[16'h50c9] <= 8'hcd;
		memory[16'h50ca] <= 8'hbc;
		memory[16'h50cb] <= 8'h5b;
		memory[16'h50cc] <= 8'h9;
		memory[16'h50cd] <= 8'h4e;
		memory[16'h50ce] <= 8'h32;
		memory[16'h50cf] <= 8'haf;
		memory[16'h50d0] <= 8'h4b;
		memory[16'h50d1] <= 8'hf2;
		memory[16'h50d2] <= 8'h5c;
		memory[16'h50d3] <= 8'h6b;
		memory[16'h50d4] <= 8'hde;
		memory[16'h50d5] <= 8'h97;
		memory[16'h50d6] <= 8'ha9;
		memory[16'h50d7] <= 8'h66;
		memory[16'h50d8] <= 8'h14;
		memory[16'h50d9] <= 8'h68;
		memory[16'h50da] <= 8'hf;
		memory[16'h50db] <= 8'h7a;
		memory[16'h50dc] <= 8'h75;
		memory[16'h50dd] <= 8'h4b;
		memory[16'h50de] <= 8'h57;
		memory[16'h50df] <= 8'hc;
		memory[16'h50e0] <= 8'hd2;
		memory[16'h50e1] <= 8'hfa;
		memory[16'h50e2] <= 8'h7c;
		memory[16'h50e3] <= 8'he4;
		memory[16'h50e4] <= 8'hf4;
		memory[16'h50e5] <= 8'h8a;
		memory[16'h50e6] <= 8'h21;
		memory[16'h50e7] <= 8'h2b;
		memory[16'h50e8] <= 8'h57;
		memory[16'h50e9] <= 8'hdd;
		memory[16'h50ea] <= 8'h86;
		memory[16'h50eb] <= 8'h60;
		memory[16'h50ec] <= 8'h2b;
		memory[16'h50ed] <= 8'hb8;
		memory[16'h50ee] <= 8'h10;
		memory[16'h50ef] <= 8'h77;
		memory[16'h50f0] <= 8'hab;
		memory[16'h50f1] <= 8'h6c;
		memory[16'h50f2] <= 8'he2;
		memory[16'h50f3] <= 8'h89;
		memory[16'h50f4] <= 8'h4;
		memory[16'h50f5] <= 8'h8c;
		memory[16'h50f6] <= 8'hef;
		memory[16'h50f7] <= 8'h18;
		memory[16'h50f8] <= 8'hf4;
		memory[16'h50f9] <= 8'hfe;
		memory[16'h50fa] <= 8'h92;
		memory[16'h50fb] <= 8'h69;
		memory[16'h50fc] <= 8'h49;
		memory[16'h50fd] <= 8'he9;
		memory[16'h50fe] <= 8'h75;
		memory[16'h50ff] <= 8'h1b;
		memory[16'h5100] <= 8'he3;
		memory[16'h5101] <= 8'hf1;
		memory[16'h5102] <= 8'h0;
		memory[16'h5103] <= 8'hd7;
		memory[16'h5104] <= 8'h7c;
		memory[16'h5105] <= 8'h21;
		memory[16'h5106] <= 8'h3;
		memory[16'h5107] <= 8'hd3;
		memory[16'h5108] <= 8'hff;
		memory[16'h5109] <= 8'h89;
		memory[16'h510a] <= 8'h34;
		memory[16'h510b] <= 8'h2a;
		memory[16'h510c] <= 8'h42;
		memory[16'h510d] <= 8'h44;
		memory[16'h510e] <= 8'ha1;
		memory[16'h510f] <= 8'hed;
		memory[16'h5110] <= 8'hb0;
		memory[16'h5111] <= 8'h84;
		memory[16'h5112] <= 8'h76;
		memory[16'h5113] <= 8'hb4;
		memory[16'h5114] <= 8'h10;
		memory[16'h5115] <= 8'h65;
		memory[16'h5116] <= 8'hcc;
		memory[16'h5117] <= 8'h4;
		memory[16'h5118] <= 8'h64;
		memory[16'h5119] <= 8'h5e;
		memory[16'h511a] <= 8'h6d;
		memory[16'h511b] <= 8'had;
		memory[16'h511c] <= 8'h47;
		memory[16'h511d] <= 8'he2;
		memory[16'h511e] <= 8'hc9;
		memory[16'h511f] <= 8'h2b;
		memory[16'h5120] <= 8'hd4;
		memory[16'h5121] <= 8'hc9;
		memory[16'h5122] <= 8'h2;
		memory[16'h5123] <= 8'h50;
		memory[16'h5124] <= 8'hea;
		memory[16'h5125] <= 8'h5;
		memory[16'h5126] <= 8'h23;
		memory[16'h5127] <= 8'he9;
		memory[16'h5128] <= 8'h8f;
		memory[16'h5129] <= 8'h57;
		memory[16'h512a] <= 8'h14;
		memory[16'h512b] <= 8'hd1;
		memory[16'h512c] <= 8'h9b;
		memory[16'h512d] <= 8'hb5;
		memory[16'h512e] <= 8'hbe;
		memory[16'h512f] <= 8'h4c;
		memory[16'h5130] <= 8'h39;
		memory[16'h5131] <= 8'h34;
		memory[16'h5132] <= 8'h0;
		memory[16'h5133] <= 8'h49;
		memory[16'h5134] <= 8'h99;
		memory[16'h5135] <= 8'hcd;
		memory[16'h5136] <= 8'h4d;
		memory[16'h5137] <= 8'hfd;
		memory[16'h5138] <= 8'h2b;
		memory[16'h5139] <= 8'hba;
		memory[16'h513a] <= 8'hab;
		memory[16'h513b] <= 8'h73;
		memory[16'h513c] <= 8'h9d;
		memory[16'h513d] <= 8'h74;
		memory[16'h513e] <= 8'h9e;
		memory[16'h513f] <= 8'h71;
		memory[16'h5140] <= 8'h3d;
		memory[16'h5141] <= 8'ha0;
		memory[16'h5142] <= 8'hc1;
		memory[16'h5143] <= 8'h27;
		memory[16'h5144] <= 8'ha6;
		memory[16'h5145] <= 8'he4;
		memory[16'h5146] <= 8'h11;
		memory[16'h5147] <= 8'h35;
		memory[16'h5148] <= 8'h3c;
		memory[16'h5149] <= 8'h25;
		memory[16'h514a] <= 8'h6;
		memory[16'h514b] <= 8'hd7;
		memory[16'h514c] <= 8'hda;
		memory[16'h514d] <= 8'hc4;
		memory[16'h514e] <= 8'h23;
		memory[16'h514f] <= 8'h14;
		memory[16'h5150] <= 8'hf8;
		memory[16'h5151] <= 8'h24;
		memory[16'h5152] <= 8'h5d;
		memory[16'h5153] <= 8'h91;
		memory[16'h5154] <= 8'hf1;
		memory[16'h5155] <= 8'hab;
		memory[16'h5156] <= 8'h8f;
		memory[16'h5157] <= 8'h1c;
		memory[16'h5158] <= 8'h65;
		memory[16'h5159] <= 8'h3a;
		memory[16'h515a] <= 8'h8f;
		memory[16'h515b] <= 8'h2;
		memory[16'h515c] <= 8'hae;
		memory[16'h515d] <= 8'h2d;
		memory[16'h515e] <= 8'h73;
		memory[16'h515f] <= 8'heb;
		memory[16'h5160] <= 8'hce;
		memory[16'h5161] <= 8'h34;
		memory[16'h5162] <= 8'h12;
		memory[16'h5163] <= 8'h74;
		memory[16'h5164] <= 8'h19;
		memory[16'h5165] <= 8'h23;
		memory[16'h5166] <= 8'ha9;
		memory[16'h5167] <= 8'h55;
		memory[16'h5168] <= 8'h48;
		memory[16'h5169] <= 8'haf;
		memory[16'h516a] <= 8'h2c;
		memory[16'h516b] <= 8'h23;
		memory[16'h516c] <= 8'h73;
		memory[16'h516d] <= 8'h50;
		memory[16'h516e] <= 8'h37;
		memory[16'h516f] <= 8'h6b;
		memory[16'h5170] <= 8'h74;
		memory[16'h5171] <= 8'h94;
		memory[16'h5172] <= 8'hfc;
		memory[16'h5173] <= 8'h65;
		memory[16'h5174] <= 8'h3f;
		memory[16'h5175] <= 8'h8b;
		memory[16'h5176] <= 8'h81;
		memory[16'h5177] <= 8'ha5;
		memory[16'h5178] <= 8'hc5;
		memory[16'h5179] <= 8'h11;
		memory[16'h517a] <= 8'ha7;
		memory[16'h517b] <= 8'h73;
		memory[16'h517c] <= 8'h3e;
		memory[16'h517d] <= 8'h1b;
		memory[16'h517e] <= 8'h5e;
		memory[16'h517f] <= 8'hc;
		memory[16'h5180] <= 8'h4f;
		memory[16'h5181] <= 8'h71;
		memory[16'h5182] <= 8'h80;
		memory[16'h5183] <= 8'h68;
		memory[16'h5184] <= 8'h94;
		memory[16'h5185] <= 8'h29;
		memory[16'h5186] <= 8'hbd;
		memory[16'h5187] <= 8'hdd;
		memory[16'h5188] <= 8'hd8;
		memory[16'h5189] <= 8'hea;
		memory[16'h518a] <= 8'h0;
		memory[16'h518b] <= 8'h4b;
		memory[16'h518c] <= 8'h3a;
		memory[16'h518d] <= 8'h37;
		memory[16'h518e] <= 8'hb6;
		memory[16'h518f] <= 8'hae;
		memory[16'h5190] <= 8'hcb;
		memory[16'h5191] <= 8'hb3;
		memory[16'h5192] <= 8'h13;
		memory[16'h5193] <= 8'hb;
		memory[16'h5194] <= 8'h3e;
		memory[16'h5195] <= 8'h94;
		memory[16'h5196] <= 8'hb0;
		memory[16'h5197] <= 8'h4;
		memory[16'h5198] <= 8'ha5;
		memory[16'h5199] <= 8'h57;
		memory[16'h519a] <= 8'h77;
		memory[16'h519b] <= 8'he4;
		memory[16'h519c] <= 8'h72;
		memory[16'h519d] <= 8'hd6;
		memory[16'h519e] <= 8'hf0;
		memory[16'h519f] <= 8'hc2;
		memory[16'h51a0] <= 8'h47;
		memory[16'h51a1] <= 8'h71;
		memory[16'h51a2] <= 8'h2a;
		memory[16'h51a3] <= 8'hdb;
		memory[16'h51a4] <= 8'h9a;
		memory[16'h51a5] <= 8'he8;
		memory[16'h51a6] <= 8'hb8;
		memory[16'h51a7] <= 8'h73;
		memory[16'h51a8] <= 8'hd2;
		memory[16'h51a9] <= 8'hb8;
		memory[16'h51aa] <= 8'hbe;
		memory[16'h51ab] <= 8'hc;
		memory[16'h51ac] <= 8'hef;
		memory[16'h51ad] <= 8'h75;
		memory[16'h51ae] <= 8'hba;
		memory[16'h51af] <= 8'hbb;
		memory[16'h51b0] <= 8'h28;
		memory[16'h51b1] <= 8'hcd;
		memory[16'h51b2] <= 8'hc6;
		memory[16'h51b3] <= 8'h66;
		memory[16'h51b4] <= 8'h61;
		memory[16'h51b5] <= 8'h76;
		memory[16'h51b6] <= 8'h6a;
		memory[16'h51b7] <= 8'h7;
		memory[16'h51b8] <= 8'hcd;
		memory[16'h51b9] <= 8'he2;
		memory[16'h51ba] <= 8'heb;
		memory[16'h51bb] <= 8'h40;
		memory[16'h51bc] <= 8'hb8;
		memory[16'h51bd] <= 8'hdb;
		memory[16'h51be] <= 8'h2;
		memory[16'h51bf] <= 8'hff;
		memory[16'h51c0] <= 8'h4c;
		memory[16'h51c1] <= 8'h2c;
		memory[16'h51c2] <= 8'hda;
		memory[16'h51c3] <= 8'he7;
		memory[16'h51c4] <= 8'h14;
		memory[16'h51c5] <= 8'h93;
		memory[16'h51c6] <= 8'h5a;
		memory[16'h51c7] <= 8'he6;
		memory[16'h51c8] <= 8'h4b;
		memory[16'h51c9] <= 8'h18;
		memory[16'h51ca] <= 8'hf2;
		memory[16'h51cb] <= 8'h3b;
		memory[16'h51cc] <= 8'h8d;
		memory[16'h51cd] <= 8'hac;
		memory[16'h51ce] <= 8'hf6;
		memory[16'h51cf] <= 8'hb5;
		memory[16'h51d0] <= 8'h79;
		memory[16'h51d1] <= 8'hbc;
		memory[16'h51d2] <= 8'h1c;
		memory[16'h51d3] <= 8'hdb;
		memory[16'h51d4] <= 8'h32;
		memory[16'h51d5] <= 8'h86;
		memory[16'h51d6] <= 8'he2;
		memory[16'h51d7] <= 8'hff;
		memory[16'h51d8] <= 8'h68;
		memory[16'h51d9] <= 8'hcd;
		memory[16'h51da] <= 8'h3f;
		memory[16'h51db] <= 8'h20;
		memory[16'h51dc] <= 8'ha8;
		memory[16'h51dd] <= 8'h41;
		memory[16'h51de] <= 8'h1f;
		memory[16'h51df] <= 8'hf5;
		memory[16'h51e0] <= 8'h6e;
		memory[16'h51e1] <= 8'hfa;
		memory[16'h51e2] <= 8'hdc;
		memory[16'h51e3] <= 8'h82;
		memory[16'h51e4] <= 8'h8d;
		memory[16'h51e5] <= 8'h36;
		memory[16'h51e6] <= 8'h69;
		memory[16'h51e7] <= 8'hd8;
		memory[16'h51e8] <= 8'h4e;
		memory[16'h51e9] <= 8'h5b;
		memory[16'h51ea] <= 8'h13;
		memory[16'h51eb] <= 8'hdc;
		memory[16'h51ec] <= 8'h8;
		memory[16'h51ed] <= 8'h9;
		memory[16'h51ee] <= 8'h91;
		memory[16'h51ef] <= 8'h81;
		memory[16'h51f0] <= 8'hc5;
		memory[16'h51f1] <= 8'had;
		memory[16'h51f2] <= 8'h5c;
		memory[16'h51f3] <= 8'hf7;
		memory[16'h51f4] <= 8'h34;
		memory[16'h51f5] <= 8'h3e;
		memory[16'h51f6] <= 8'hf7;
		memory[16'h51f7] <= 8'h9c;
		memory[16'h51f8] <= 8'hb;
		memory[16'h51f9] <= 8'h36;
		memory[16'h51fa] <= 8'hbd;
		memory[16'h51fb] <= 8'hb4;
		memory[16'h51fc] <= 8'h78;
		memory[16'h51fd] <= 8'hdc;
		memory[16'h51fe] <= 8'ha9;
		memory[16'h51ff] <= 8'he6;
		memory[16'h5200] <= 8'hd6;
		memory[16'h5201] <= 8'h85;
		memory[16'h5202] <= 8'h68;
		memory[16'h5203] <= 8'h63;
		memory[16'h5204] <= 8'hbb;
		memory[16'h5205] <= 8'hd1;
		memory[16'h5206] <= 8'h3c;
		memory[16'h5207] <= 8'h9;
		memory[16'h5208] <= 8'h2d;
		memory[16'h5209] <= 8'h4f;
		memory[16'h520a] <= 8'he5;
		memory[16'h520b] <= 8'h35;
		memory[16'h520c] <= 8'h59;
		memory[16'h520d] <= 8'h77;
		memory[16'h520e] <= 8'hb6;
		memory[16'h520f] <= 8'h1e;
		memory[16'h5210] <= 8'h24;
		memory[16'h5211] <= 8'h13;
		memory[16'h5212] <= 8'h16;
		memory[16'h5213] <= 8'h58;
		memory[16'h5214] <= 8'h51;
		memory[16'h5215] <= 8'hd;
		memory[16'h5216] <= 8'hf5;
		memory[16'h5217] <= 8'h5d;
		memory[16'h5218] <= 8'h43;
		memory[16'h5219] <= 8'hb2;
		memory[16'h521a] <= 8'h11;
		memory[16'h521b] <= 8'hbb;
		memory[16'h521c] <= 8'h8e;
		memory[16'h521d] <= 8'hba;
		memory[16'h521e] <= 8'ha1;
		memory[16'h521f] <= 8'h65;
		memory[16'h5220] <= 8'h3f;
		memory[16'h5221] <= 8'ha;
		memory[16'h5222] <= 8'hc8;
		memory[16'h5223] <= 8'hfa;
		memory[16'h5224] <= 8'hdb;
		memory[16'h5225] <= 8'h4;
		memory[16'h5226] <= 8'h3;
		memory[16'h5227] <= 8'h8;
		memory[16'h5228] <= 8'h54;
		memory[16'h5229] <= 8'he9;
		memory[16'h522a] <= 8'h3d;
		memory[16'h522b] <= 8'had;
		memory[16'h522c] <= 8'h60;
		memory[16'h522d] <= 8'hf4;
		memory[16'h522e] <= 8'hcb;
		memory[16'h522f] <= 8'h84;
		memory[16'h5230] <= 8'h7;
		memory[16'h5231] <= 8'he1;
		memory[16'h5232] <= 8'hdd;
		memory[16'h5233] <= 8'h58;
		memory[16'h5234] <= 8'hee;
		memory[16'h5235] <= 8'hd2;
		memory[16'h5236] <= 8'hb5;
		memory[16'h5237] <= 8'h32;
		memory[16'h5238] <= 8'h84;
		memory[16'h5239] <= 8'hc6;
		memory[16'h523a] <= 8'hed;
		memory[16'h523b] <= 8'h12;
		memory[16'h523c] <= 8'h80;
		memory[16'h523d] <= 8'h8f;
		memory[16'h523e] <= 8'h77;
		memory[16'h523f] <= 8'hbf;
		memory[16'h5240] <= 8'h99;
		memory[16'h5241] <= 8'h40;
		memory[16'h5242] <= 8'hb9;
		memory[16'h5243] <= 8'h74;
		memory[16'h5244] <= 8'h44;
		memory[16'h5245] <= 8'hbd;
		memory[16'h5246] <= 8'h7d;
		memory[16'h5247] <= 8'h98;
		memory[16'h5248] <= 8'ha6;
		memory[16'h5249] <= 8'hba;
		memory[16'h524a] <= 8'h45;
		memory[16'h524b] <= 8'h6;
		memory[16'h524c] <= 8'hae;
		memory[16'h524d] <= 8'h11;
		memory[16'h524e] <= 8'h8a;
		memory[16'h524f] <= 8'hb5;
		memory[16'h5250] <= 8'hf2;
		memory[16'h5251] <= 8'h67;
		memory[16'h5252] <= 8'he;
		memory[16'h5253] <= 8'he1;
		memory[16'h5254] <= 8'h39;
		memory[16'h5255] <= 8'hc3;
		memory[16'h5256] <= 8'h13;
		memory[16'h5257] <= 8'hbd;
		memory[16'h5258] <= 8'h8a;
		memory[16'h5259] <= 8'h0;
		memory[16'h525a] <= 8'hd0;
		memory[16'h525b] <= 8'ha;
		memory[16'h525c] <= 8'h8f;
		memory[16'h525d] <= 8'h47;
		memory[16'h525e] <= 8'hca;
		memory[16'h525f] <= 8'h28;
		memory[16'h5260] <= 8'h87;
		memory[16'h5261] <= 8'h83;
		memory[16'h5262] <= 8'h9d;
		memory[16'h5263] <= 8'hcc;
		memory[16'h5264] <= 8'h40;
		memory[16'h5265] <= 8'h1a;
		memory[16'h5266] <= 8'h64;
		memory[16'h5267] <= 8'he6;
		memory[16'h5268] <= 8'hd4;
		memory[16'h5269] <= 8'haa;
		memory[16'h526a] <= 8'hec;
		memory[16'h526b] <= 8'h83;
		memory[16'h526c] <= 8'hbb;
		memory[16'h526d] <= 8'h77;
		memory[16'h526e] <= 8'h38;
		memory[16'h526f] <= 8'had;
		memory[16'h5270] <= 8'hde;
		memory[16'h5271] <= 8'h46;
		memory[16'h5272] <= 8'h8e;
		memory[16'h5273] <= 8'h18;
		memory[16'h5274] <= 8'ha;
		memory[16'h5275] <= 8'ha1;
		memory[16'h5276] <= 8'hd5;
		memory[16'h5277] <= 8'h94;
		memory[16'h5278] <= 8'ha2;
		memory[16'h5279] <= 8'ha5;
		memory[16'h527a] <= 8'h9e;
		memory[16'h527b] <= 8'h31;
		memory[16'h527c] <= 8'hed;
		memory[16'h527d] <= 8'h68;
		memory[16'h527e] <= 8'h5a;
		memory[16'h527f] <= 8'h74;
		memory[16'h5280] <= 8'hec;
		memory[16'h5281] <= 8'hf7;
		memory[16'h5282] <= 8'h40;
		memory[16'h5283] <= 8'h2c;
		memory[16'h5284] <= 8'h11;
		memory[16'h5285] <= 8'ha5;
		memory[16'h5286] <= 8'h13;
		memory[16'h5287] <= 8'he5;
		memory[16'h5288] <= 8'h4f;
		memory[16'h5289] <= 8'hff;
		memory[16'h528a] <= 8'h68;
		memory[16'h528b] <= 8'ha;
		memory[16'h528c] <= 8'h76;
		memory[16'h528d] <= 8'ha1;
		memory[16'h528e] <= 8'hb7;
		memory[16'h528f] <= 8'h55;
		memory[16'h5290] <= 8'he7;
		memory[16'h5291] <= 8'h46;
		memory[16'h5292] <= 8'h6d;
		memory[16'h5293] <= 8'hf1;
		memory[16'h5294] <= 8'he7;
		memory[16'h5295] <= 8'h42;
		memory[16'h5296] <= 8'h85;
		memory[16'h5297] <= 8'h89;
		memory[16'h5298] <= 8'he8;
		memory[16'h5299] <= 8'h24;
		memory[16'h529a] <= 8'hbb;
		memory[16'h529b] <= 8'hd5;
		memory[16'h529c] <= 8'h8c;
		memory[16'h529d] <= 8'h15;
		memory[16'h529e] <= 8'h49;
		memory[16'h529f] <= 8'h78;
		memory[16'h52a0] <= 8'hc;
		memory[16'h52a1] <= 8'h8a;
		memory[16'h52a2] <= 8'ha5;
		memory[16'h52a3] <= 8'h1d;
		memory[16'h52a4] <= 8'h2f;
		memory[16'h52a5] <= 8'hb8;
		memory[16'h52a6] <= 8'h2;
		memory[16'h52a7] <= 8'h7e;
		memory[16'h52a8] <= 8'hb7;
		memory[16'h52a9] <= 8'h6b;
		memory[16'h52aa] <= 8'h88;
		memory[16'h52ab] <= 8'h2e;
		memory[16'h52ac] <= 8'hc;
		memory[16'h52ad] <= 8'h3f;
		memory[16'h52ae] <= 8'h83;
		memory[16'h52af] <= 8'hf3;
		memory[16'h52b0] <= 8'h85;
		memory[16'h52b1] <= 8'hf0;
		memory[16'h52b2] <= 8'he5;
		memory[16'h52b3] <= 8'h6d;
		memory[16'h52b4] <= 8'h32;
		memory[16'h52b5] <= 8'h6a;
		memory[16'h52b6] <= 8'hf6;
		memory[16'h52b7] <= 8'h1a;
		memory[16'h52b8] <= 8'h8e;
		memory[16'h52b9] <= 8'hb1;
		memory[16'h52ba] <= 8'hef;
		memory[16'h52bb] <= 8'h1b;
		memory[16'h52bc] <= 8'hc6;
		memory[16'h52bd] <= 8'h39;
		memory[16'h52be] <= 8'h93;
		memory[16'h52bf] <= 8'hd2;
		memory[16'h52c0] <= 8'hc3;
		memory[16'h52c1] <= 8'h38;
		memory[16'h52c2] <= 8'hef;
		memory[16'h52c3] <= 8'hf2;
		memory[16'h52c4] <= 8'hf0;
		memory[16'h52c5] <= 8'hf2;
		memory[16'h52c6] <= 8'h70;
		memory[16'h52c7] <= 8'ha8;
		memory[16'h52c8] <= 8'h5d;
		memory[16'h52c9] <= 8'hf8;
		memory[16'h52ca] <= 8'hd6;
		memory[16'h52cb] <= 8'h69;
		memory[16'h52cc] <= 8'h37;
		memory[16'h52cd] <= 8'h59;
		memory[16'h52ce] <= 8'h5c;
		memory[16'h52cf] <= 8'hbd;
		memory[16'h52d0] <= 8'h49;
		memory[16'h52d1] <= 8'h41;
		memory[16'h52d2] <= 8'h2a;
		memory[16'h52d3] <= 8'h7b;
		memory[16'h52d4] <= 8'hac;
		memory[16'h52d5] <= 8'h20;
		memory[16'h52d6] <= 8'h96;
		memory[16'h52d7] <= 8'h3a;
		memory[16'h52d8] <= 8'hd2;
		memory[16'h52d9] <= 8'h85;
		memory[16'h52da] <= 8'h55;
		memory[16'h52db] <= 8'h98;
		memory[16'h52dc] <= 8'hbe;
		memory[16'h52dd] <= 8'he9;
		memory[16'h52de] <= 8'h6b;
		memory[16'h52df] <= 8'h81;
		memory[16'h52e0] <= 8'h21;
		memory[16'h52e1] <= 8'h5a;
		memory[16'h52e2] <= 8'h73;
		memory[16'h52e3] <= 8'h12;
		memory[16'h52e4] <= 8'h4c;
		memory[16'h52e5] <= 8'he3;
		memory[16'h52e6] <= 8'hba;
		memory[16'h52e7] <= 8'ha9;
		memory[16'h52e8] <= 8'hdb;
		memory[16'h52e9] <= 8'h90;
		memory[16'h52ea] <= 8'h12;
		memory[16'h52eb] <= 8'h13;
		memory[16'h52ec] <= 8'he9;
		memory[16'h52ed] <= 8'h6f;
		memory[16'h52ee] <= 8'hd0;
		memory[16'h52ef] <= 8'h32;
		memory[16'h52f0] <= 8'hb0;
		memory[16'h52f1] <= 8'hfa;
		memory[16'h52f2] <= 8'had;
		memory[16'h52f3] <= 8'h5c;
		memory[16'h52f4] <= 8'h1a;
		memory[16'h52f5] <= 8'h43;
		memory[16'h52f6] <= 8'h97;
		memory[16'h52f7] <= 8'hec;
		memory[16'h52f8] <= 8'hc9;
		memory[16'h52f9] <= 8'hec;
		memory[16'h52fa] <= 8'h85;
		memory[16'h52fb] <= 8'h87;
		memory[16'h52fc] <= 8'hd5;
		memory[16'h52fd] <= 8'hf0;
		memory[16'h52fe] <= 8'h9;
		memory[16'h52ff] <= 8'hf7;
		memory[16'h5300] <= 8'h4a;
		memory[16'h5301] <= 8'h7c;
		memory[16'h5302] <= 8'h9;
		memory[16'h5303] <= 8'h97;
		memory[16'h5304] <= 8'h60;
		memory[16'h5305] <= 8'hc3;
		memory[16'h5306] <= 8'h40;
		memory[16'h5307] <= 8'h3b;
		memory[16'h5308] <= 8'h53;
		memory[16'h5309] <= 8'h53;
		memory[16'h530a] <= 8'h4e;
		memory[16'h530b] <= 8'h3c;
		memory[16'h530c] <= 8'hc2;
		memory[16'h530d] <= 8'h1e;
		memory[16'h530e] <= 8'h6e;
		memory[16'h530f] <= 8'h72;
		memory[16'h5310] <= 8'h18;
		memory[16'h5311] <= 8'h1b;
		memory[16'h5312] <= 8'hcf;
		memory[16'h5313] <= 8'h33;
		memory[16'h5314] <= 8'h5f;
		memory[16'h5315] <= 8'h66;
		memory[16'h5316] <= 8'h1f;
		memory[16'h5317] <= 8'h28;
		memory[16'h5318] <= 8'h52;
		memory[16'h5319] <= 8'ha4;
		memory[16'h531a] <= 8'haf;
		memory[16'h531b] <= 8'h28;
		memory[16'h531c] <= 8'h94;
		memory[16'h531d] <= 8'hb8;
		memory[16'h531e] <= 8'h1f;
		memory[16'h531f] <= 8'hdf;
		memory[16'h5320] <= 8'h35;
		memory[16'h5321] <= 8'h28;
		memory[16'h5322] <= 8'h76;
		memory[16'h5323] <= 8'h95;
		memory[16'h5324] <= 8'heb;
		memory[16'h5325] <= 8'hb6;
		memory[16'h5326] <= 8'hd0;
		memory[16'h5327] <= 8'h3e;
		memory[16'h5328] <= 8'h9;
		memory[16'h5329] <= 8'h1f;
		memory[16'h532a] <= 8'h7a;
		memory[16'h532b] <= 8'hcb;
		memory[16'h532c] <= 8'h3d;
		memory[16'h532d] <= 8'he8;
		memory[16'h532e] <= 8'h3e;
		memory[16'h532f] <= 8'h56;
		memory[16'h5330] <= 8'h3;
		memory[16'h5331] <= 8'hd;
		memory[16'h5332] <= 8'h89;
		memory[16'h5333] <= 8'h62;
		memory[16'h5334] <= 8'h73;
		memory[16'h5335] <= 8'ha8;
		memory[16'h5336] <= 8'h8a;
		memory[16'h5337] <= 8'hc5;
		memory[16'h5338] <= 8'h4d;
		memory[16'h5339] <= 8'h3a;
		memory[16'h533a] <= 8'hed;
		memory[16'h533b] <= 8'he1;
		memory[16'h533c] <= 8'hf2;
		memory[16'h533d] <= 8'hc;
		memory[16'h533e] <= 8'hc0;
		memory[16'h533f] <= 8'h27;
		memory[16'h5340] <= 8'h34;
		memory[16'h5341] <= 8'h36;
		memory[16'h5342] <= 8'hbc;
		memory[16'h5343] <= 8'h1f;
		memory[16'h5344] <= 8'hed;
		memory[16'h5345] <= 8'h8d;
		memory[16'h5346] <= 8'h5d;
		memory[16'h5347] <= 8'hf6;
		memory[16'h5348] <= 8'hac;
		memory[16'h5349] <= 8'hd7;
		memory[16'h534a] <= 8'hc2;
		memory[16'h534b] <= 8'he9;
		memory[16'h534c] <= 8'hbf;
		memory[16'h534d] <= 8'h0;
		memory[16'h534e] <= 8'h3f;
		memory[16'h534f] <= 8'hc3;
		memory[16'h5350] <= 8'hd;
		memory[16'h5351] <= 8'hc8;
		memory[16'h5352] <= 8'h25;
		memory[16'h5353] <= 8'h80;
		memory[16'h5354] <= 8'h71;
		memory[16'h5355] <= 8'hb0;
		memory[16'h5356] <= 8'h45;
		memory[16'h5357] <= 8'hbe;
		memory[16'h5358] <= 8'hea;
		memory[16'h5359] <= 8'h33;
		memory[16'h535a] <= 8'h9f;
		memory[16'h535b] <= 8'hdc;
		memory[16'h535c] <= 8'h3f;
		memory[16'h535d] <= 8'h60;
		memory[16'h535e] <= 8'h4;
		memory[16'h535f] <= 8'h74;
		memory[16'h5360] <= 8'h96;
		memory[16'h5361] <= 8'hc0;
		memory[16'h5362] <= 8'h93;
		memory[16'h5363] <= 8'h83;
		memory[16'h5364] <= 8'h4d;
		memory[16'h5365] <= 8'hf1;
		memory[16'h5366] <= 8'h7a;
		memory[16'h5367] <= 8'hf9;
		memory[16'h5368] <= 8'hc8;
		memory[16'h5369] <= 8'h3c;
		memory[16'h536a] <= 8'he3;
		memory[16'h536b] <= 8'h88;
		memory[16'h536c] <= 8'h3c;
		memory[16'h536d] <= 8'h22;
		memory[16'h536e] <= 8'h4b;
		memory[16'h536f] <= 8'h49;
		memory[16'h5370] <= 8'heb;
		memory[16'h5371] <= 8'h70;
		memory[16'h5372] <= 8'hc9;
		memory[16'h5373] <= 8'h5c;
		memory[16'h5374] <= 8'h20;
		memory[16'h5375] <= 8'he;
		memory[16'h5376] <= 8'h1a;
		memory[16'h5377] <= 8'ha;
		memory[16'h5378] <= 8'h41;
		memory[16'h5379] <= 8'hb9;
		memory[16'h537a] <= 8'he7;
		memory[16'h537b] <= 8'h81;
		memory[16'h537c] <= 8'h19;
		memory[16'h537d] <= 8'heb;
		memory[16'h537e] <= 8'hf5;
		memory[16'h537f] <= 8'hb0;
		memory[16'h5380] <= 8'hab;
		memory[16'h5381] <= 8'h88;
		memory[16'h5382] <= 8'h33;
		memory[16'h5383] <= 8'hf9;
		memory[16'h5384] <= 8'h79;
		memory[16'h5385] <= 8'had;
		memory[16'h5386] <= 8'hf2;
		memory[16'h5387] <= 8'h42;
		memory[16'h5388] <= 8'he9;
		memory[16'h5389] <= 8'hd5;
		memory[16'h538a] <= 8'hca;
		memory[16'h538b] <= 8'h25;
		memory[16'h538c] <= 8'hf8;
		memory[16'h538d] <= 8'h15;
		memory[16'h538e] <= 8'h6e;
		memory[16'h538f] <= 8'he3;
		memory[16'h5390] <= 8'h85;
		memory[16'h5391] <= 8'h37;
		memory[16'h5392] <= 8'h3f;
		memory[16'h5393] <= 8'ha6;
		memory[16'h5394] <= 8'h46;
		memory[16'h5395] <= 8'h59;
		memory[16'h5396] <= 8'hb0;
		memory[16'h5397] <= 8'h87;
		memory[16'h5398] <= 8'h12;
		memory[16'h5399] <= 8'h97;
		memory[16'h539a] <= 8'h8;
		memory[16'h539b] <= 8'h2c;
		memory[16'h539c] <= 8'h82;
		memory[16'h539d] <= 8'hfd;
		memory[16'h539e] <= 8'hdc;
		memory[16'h539f] <= 8'h2e;
		memory[16'h53a0] <= 8'h86;
		memory[16'h53a1] <= 8'hf;
		memory[16'h53a2] <= 8'h27;
		memory[16'h53a3] <= 8'hff;
		memory[16'h53a4] <= 8'hbd;
		memory[16'h53a5] <= 8'h19;
		memory[16'h53a6] <= 8'h41;
		memory[16'h53a7] <= 8'ha6;
		memory[16'h53a8] <= 8'hef;
		memory[16'h53a9] <= 8'hb;
		memory[16'h53aa] <= 8'hcc;
		memory[16'h53ab] <= 8'he7;
		memory[16'h53ac] <= 8'h20;
		memory[16'h53ad] <= 8'h3a;
		memory[16'h53ae] <= 8'hca;
		memory[16'h53af] <= 8'ha6;
		memory[16'h53b0] <= 8'h72;
		memory[16'h53b1] <= 8'h9;
		memory[16'h53b2] <= 8'h4c;
		memory[16'h53b3] <= 8'hb8;
		memory[16'h53b4] <= 8'h62;
		memory[16'h53b5] <= 8'hfc;
		memory[16'h53b6] <= 8'h3f;
		memory[16'h53b7] <= 8'h74;
		memory[16'h53b8] <= 8'h94;
		memory[16'h53b9] <= 8'h48;
		memory[16'h53ba] <= 8'ha0;
		memory[16'h53bb] <= 8'h16;
		memory[16'h53bc] <= 8'h45;
		memory[16'h53bd] <= 8'h7c;
		memory[16'h53be] <= 8'h44;
		memory[16'h53bf] <= 8'hcb;
		memory[16'h53c0] <= 8'h8c;
		memory[16'h53c1] <= 8'h6b;
		memory[16'h53c2] <= 8'hcb;
		memory[16'h53c3] <= 8'h49;
		memory[16'h53c4] <= 8'h85;
		memory[16'h53c5] <= 8'hc;
		memory[16'h53c6] <= 8'hef;
		memory[16'h53c7] <= 8'h74;
		memory[16'h53c8] <= 8'h18;
		memory[16'h53c9] <= 8'hbb;
		memory[16'h53ca] <= 8'h5b;
		memory[16'h53cb] <= 8'h38;
		memory[16'h53cc] <= 8'hf6;
		memory[16'h53cd] <= 8'h25;
		memory[16'h53ce] <= 8'hde;
		memory[16'h53cf] <= 8'h68;
		memory[16'h53d0] <= 8'h2e;
		memory[16'h53d1] <= 8'h2a;
		memory[16'h53d2] <= 8'h20;
		memory[16'h53d3] <= 8'h90;
		memory[16'h53d4] <= 8'h27;
		memory[16'h53d5] <= 8'h5f;
		memory[16'h53d6] <= 8'h4;
		memory[16'h53d7] <= 8'hbb;
		memory[16'h53d8] <= 8'ha7;
		memory[16'h53d9] <= 8'ha5;
		memory[16'h53da] <= 8'hd1;
		memory[16'h53db] <= 8'hed;
		memory[16'h53dc] <= 8'h21;
		memory[16'h53dd] <= 8'h16;
		memory[16'h53de] <= 8'hb8;
		memory[16'h53df] <= 8'had;
		memory[16'h53e0] <= 8'h81;
		memory[16'h53e1] <= 8'h83;
		memory[16'h53e2] <= 8'hf6;
		memory[16'h53e3] <= 8'h6;
		memory[16'h53e4] <= 8'h90;
		memory[16'h53e5] <= 8'he6;
		memory[16'h53e6] <= 8'h7a;
		memory[16'h53e7] <= 8'ha8;
		memory[16'h53e8] <= 8'ha1;
		memory[16'h53e9] <= 8'hd5;
		memory[16'h53ea] <= 8'he0;
		memory[16'h53eb] <= 8'h97;
		memory[16'h53ec] <= 8'hfa;
		memory[16'h53ed] <= 8'hbf;
		memory[16'h53ee] <= 8'hff;
		memory[16'h53ef] <= 8'h28;
		memory[16'h53f0] <= 8'he9;
		memory[16'h53f1] <= 8'h1f;
		memory[16'h53f2] <= 8'hb8;
		memory[16'h53f3] <= 8'h10;
		memory[16'h53f4] <= 8'h7f;
		memory[16'h53f5] <= 8'hbd;
		memory[16'h53f6] <= 8'hcb;
		memory[16'h53f7] <= 8'h26;
		memory[16'h53f8] <= 8'h62;
		memory[16'h53f9] <= 8'h9d;
		memory[16'h53fa] <= 8'h13;
		memory[16'h53fb] <= 8'h83;
		memory[16'h53fc] <= 8'hb3;
		memory[16'h53fd] <= 8'hcc;
		memory[16'h53fe] <= 8'h31;
		memory[16'h53ff] <= 8'h34;
		memory[16'h5400] <= 8'h4f;
		memory[16'h5401] <= 8'h27;
		memory[16'h5402] <= 8'h3b;
		memory[16'h5403] <= 8'hdf;
		memory[16'h5404] <= 8'hd;
		memory[16'h5405] <= 8'hb5;
		memory[16'h5406] <= 8'h87;
		memory[16'h5407] <= 8'haf;
		memory[16'h5408] <= 8'h8b;
		memory[16'h5409] <= 8'h68;
		memory[16'h540a] <= 8'h46;
		memory[16'h540b] <= 8'h85;
		memory[16'h540c] <= 8'h27;
		memory[16'h540d] <= 8'h46;
		memory[16'h540e] <= 8'hae;
		memory[16'h540f] <= 8'h10;
		memory[16'h5410] <= 8'h65;
		memory[16'h5411] <= 8'h66;
		memory[16'h5412] <= 8'h21;
		memory[16'h5413] <= 8'he4;
		memory[16'h5414] <= 8'h23;
		memory[16'h5415] <= 8'hec;
		memory[16'h5416] <= 8'hb;
		memory[16'h5417] <= 8'h85;
		memory[16'h5418] <= 8'h89;
		memory[16'h5419] <= 8'h1e;
		memory[16'h541a] <= 8'h9;
		memory[16'h541b] <= 8'h3c;
		memory[16'h541c] <= 8'hea;
		memory[16'h541d] <= 8'h3a;
		memory[16'h541e] <= 8'h71;
		memory[16'h541f] <= 8'h3a;
		memory[16'h5420] <= 8'h61;
		memory[16'h5421] <= 8'hac;
		memory[16'h5422] <= 8'h19;
		memory[16'h5423] <= 8'h6f;
		memory[16'h5424] <= 8'h61;
		memory[16'h5425] <= 8'ha1;
		memory[16'h5426] <= 8'h1e;
		memory[16'h5427] <= 8'hec;
		memory[16'h5428] <= 8'h9;
		memory[16'h5429] <= 8'h64;
		memory[16'h542a] <= 8'h72;
		memory[16'h542b] <= 8'h30;
		memory[16'h542c] <= 8'haa;
		memory[16'h542d] <= 8'h20;
		memory[16'h542e] <= 8'h40;
		memory[16'h542f] <= 8'h10;
		memory[16'h5430] <= 8'h86;
		memory[16'h5431] <= 8'h61;
		memory[16'h5432] <= 8'hf4;
		memory[16'h5433] <= 8'haa;
		memory[16'h5434] <= 8'h4e;
		memory[16'h5435] <= 8'hff;
		memory[16'h5436] <= 8'h2f;
		memory[16'h5437] <= 8'hd7;
		memory[16'h5438] <= 8'h1e;
		memory[16'h5439] <= 8'h38;
		memory[16'h543a] <= 8'h14;
		memory[16'h543b] <= 8'h8;
		memory[16'h543c] <= 8'h72;
		memory[16'h543d] <= 8'h85;
		memory[16'h543e] <= 8'h42;
		memory[16'h543f] <= 8'hd4;
		memory[16'h5440] <= 8'h31;
		memory[16'h5441] <= 8'h5c;
		memory[16'h5442] <= 8'h43;
		memory[16'h5443] <= 8'h92;
		memory[16'h5444] <= 8'hfd;
		memory[16'h5445] <= 8'h61;
		memory[16'h5446] <= 8'h7f;
		memory[16'h5447] <= 8'h6;
		memory[16'h5448] <= 8'hc5;
		memory[16'h5449] <= 8'hf1;
		memory[16'h544a] <= 8'h36;
		memory[16'h544b] <= 8'h70;
		memory[16'h544c] <= 8'h11;
		memory[16'h544d] <= 8'h76;
		memory[16'h544e] <= 8'h80;
		memory[16'h544f] <= 8'h97;
		memory[16'h5450] <= 8'hd8;
		memory[16'h5451] <= 8'h74;
		memory[16'h5452] <= 8'h41;
		memory[16'h5453] <= 8'h26;
		memory[16'h5454] <= 8'h74;
		memory[16'h5455] <= 8'h71;
		memory[16'h5456] <= 8'hfd;
		memory[16'h5457] <= 8'h92;
		memory[16'h5458] <= 8'ha9;
		memory[16'h5459] <= 8'h11;
		memory[16'h545a] <= 8'h9a;
		memory[16'h545b] <= 8'h1c;
		memory[16'h545c] <= 8'h96;
		memory[16'h545d] <= 8'hdd;
		memory[16'h545e] <= 8'hf0;
		memory[16'h545f] <= 8'hc7;
		memory[16'h5460] <= 8'h39;
		memory[16'h5461] <= 8'h33;
		memory[16'h5462] <= 8'h5a;
		memory[16'h5463] <= 8'h36;
		memory[16'h5464] <= 8'h94;
		memory[16'h5465] <= 8'hd9;
		memory[16'h5466] <= 8'h3c;
		memory[16'h5467] <= 8'h59;
		memory[16'h5468] <= 8'hca;
		memory[16'h5469] <= 8'h72;
		memory[16'h546a] <= 8'hc9;
		memory[16'h546b] <= 8'hdb;
		memory[16'h546c] <= 8'he8;
		memory[16'h546d] <= 8'h49;
		memory[16'h546e] <= 8'h72;
		memory[16'h546f] <= 8'hc0;
		memory[16'h5470] <= 8'hbe;
		memory[16'h5471] <= 8'hb4;
		memory[16'h5472] <= 8'he6;
		memory[16'h5473] <= 8'h32;
		memory[16'h5474] <= 8'h25;
		memory[16'h5475] <= 8'he4;
		memory[16'h5476] <= 8'hc4;
		memory[16'h5477] <= 8'hce;
		memory[16'h5478] <= 8'hf5;
		memory[16'h5479] <= 8'h5e;
		memory[16'h547a] <= 8'hea;
		memory[16'h547b] <= 8'h8c;
		memory[16'h547c] <= 8'h3b;
		memory[16'h547d] <= 8'hda;
		memory[16'h547e] <= 8'h53;
		memory[16'h547f] <= 8'h74;
		memory[16'h5480] <= 8'hd;
		memory[16'h5481] <= 8'had;
		memory[16'h5482] <= 8'haa;
		memory[16'h5483] <= 8'ha1;
		memory[16'h5484] <= 8'h86;
		memory[16'h5485] <= 8'he6;
		memory[16'h5486] <= 8'hfb;
		memory[16'h5487] <= 8'h50;
		memory[16'h5488] <= 8'h58;
		memory[16'h5489] <= 8'hc4;
		memory[16'h548a] <= 8'h2b;
		memory[16'h548b] <= 8'h41;
		memory[16'h548c] <= 8'he;
		memory[16'h548d] <= 8'h9e;
		memory[16'h548e] <= 8'h1;
		memory[16'h548f] <= 8'hcc;
		memory[16'h5490] <= 8'h52;
		memory[16'h5491] <= 8'he8;
		memory[16'h5492] <= 8'hfe;
		memory[16'h5493] <= 8'h77;
		memory[16'h5494] <= 8'hcc;
		memory[16'h5495] <= 8'hc2;
		memory[16'h5496] <= 8'h45;
		memory[16'h5497] <= 8'hc1;
		memory[16'h5498] <= 8'h20;
		memory[16'h5499] <= 8'h30;
		memory[16'h549a] <= 8'h4d;
		memory[16'h549b] <= 8'h5c;
		memory[16'h549c] <= 8'ha;
		memory[16'h549d] <= 8'ha1;
		memory[16'h549e] <= 8'hd0;
		memory[16'h549f] <= 8'h18;
		memory[16'h54a0] <= 8'h4e;
		memory[16'h54a1] <= 8'h7b;
		memory[16'h54a2] <= 8'hb9;
		memory[16'h54a3] <= 8'hd5;
		memory[16'h54a4] <= 8'h61;
		memory[16'h54a5] <= 8'hb4;
		memory[16'h54a6] <= 8'h25;
		memory[16'h54a7] <= 8'hba;
		memory[16'h54a8] <= 8'h79;
		memory[16'h54a9] <= 8'h51;
		memory[16'h54aa] <= 8'hfb;
		memory[16'h54ab] <= 8'h87;
		memory[16'h54ac] <= 8'hef;
		memory[16'h54ad] <= 8'hfc;
		memory[16'h54ae] <= 8'h53;
		memory[16'h54af] <= 8'h41;
		memory[16'h54b0] <= 8'he4;
		memory[16'h54b1] <= 8'h51;
		memory[16'h54b2] <= 8'hb8;
		memory[16'h54b3] <= 8'hb0;
		memory[16'h54b4] <= 8'h13;
		memory[16'h54b5] <= 8'hfd;
		memory[16'h54b6] <= 8'h72;
		memory[16'h54b7] <= 8'h33;
		memory[16'h54b8] <= 8'h2d;
		memory[16'h54b9] <= 8'hbf;
		memory[16'h54ba] <= 8'h8f;
		memory[16'h54bb] <= 8'h38;
		memory[16'h54bc] <= 8'h60;
		memory[16'h54bd] <= 8'h60;
		memory[16'h54be] <= 8'h50;
		memory[16'h54bf] <= 8'haf;
		memory[16'h54c0] <= 8'hdb;
		memory[16'h54c1] <= 8'h9;
		memory[16'h54c2] <= 8'h84;
		memory[16'h54c3] <= 8'h3c;
		memory[16'h54c4] <= 8'hbe;
		memory[16'h54c5] <= 8'ha9;
		memory[16'h54c6] <= 8'hf6;
		memory[16'h54c7] <= 8'h37;
		memory[16'h54c8] <= 8'hfa;
		memory[16'h54c9] <= 8'hf1;
		memory[16'h54ca] <= 8'hbe;
		memory[16'h54cb] <= 8'he9;
		memory[16'h54cc] <= 8'hee;
		memory[16'h54cd] <= 8'h11;
		memory[16'h54ce] <= 8'h2a;
		memory[16'h54cf] <= 8'hd2;
		memory[16'h54d0] <= 8'h62;
		memory[16'h54d1] <= 8'he2;
		memory[16'h54d2] <= 8'h83;
		memory[16'h54d3] <= 8'h75;
		memory[16'h54d4] <= 8'he0;
		memory[16'h54d5] <= 8'hf5;
		memory[16'h54d6] <= 8'ha8;
		memory[16'h54d7] <= 8'hd;
		memory[16'h54d8] <= 8'hb4;
		memory[16'h54d9] <= 8'h38;
		memory[16'h54da] <= 8'h45;
		memory[16'h54db] <= 8'h15;
		memory[16'h54dc] <= 8'h98;
		memory[16'h54dd] <= 8'h95;
		memory[16'h54de] <= 8'hc4;
		memory[16'h54df] <= 8'h73;
		memory[16'h54e0] <= 8'h9f;
		memory[16'h54e1] <= 8'h48;
		memory[16'h54e2] <= 8'haf;
		memory[16'h54e3] <= 8'h5d;
		memory[16'h54e4] <= 8'hf1;
		memory[16'h54e5] <= 8'ha6;
		memory[16'h54e6] <= 8'h94;
		memory[16'h54e7] <= 8'hec;
		memory[16'h54e8] <= 8'h97;
		memory[16'h54e9] <= 8'h52;
		memory[16'h54ea] <= 8'hd5;
		memory[16'h54eb] <= 8'h85;
		memory[16'h54ec] <= 8'h63;
		memory[16'h54ed] <= 8'h0;
		memory[16'h54ee] <= 8'h58;
		memory[16'h54ef] <= 8'hc5;
		memory[16'h54f0] <= 8'he2;
		memory[16'h54f1] <= 8'hdb;
		memory[16'h54f2] <= 8'h3a;
		memory[16'h54f3] <= 8'hc2;
		memory[16'h54f4] <= 8'hd0;
		memory[16'h54f5] <= 8'he2;
		memory[16'h54f6] <= 8'hd0;
		memory[16'h54f7] <= 8'h84;
		memory[16'h54f8] <= 8'h1a;
		memory[16'h54f9] <= 8'h15;
		memory[16'h54fa] <= 8'h99;
		memory[16'h54fb] <= 8'hb2;
		memory[16'h54fc] <= 8'hab;
		memory[16'h54fd] <= 8'h5d;
		memory[16'h54fe] <= 8'h25;
		memory[16'h54ff] <= 8'h4a;
		memory[16'h5500] <= 8'ha5;
		memory[16'h5501] <= 8'hd5;
		memory[16'h5502] <= 8'ha7;
		memory[16'h5503] <= 8'h97;
		memory[16'h5504] <= 8'h7b;
		memory[16'h5505] <= 8'h3b;
		memory[16'h5506] <= 8'h83;
		memory[16'h5507] <= 8'h12;
		memory[16'h5508] <= 8'h8d;
		memory[16'h5509] <= 8'h58;
		memory[16'h550a] <= 8'h98;
		memory[16'h550b] <= 8'hf0;
		memory[16'h550c] <= 8'h58;
		memory[16'h550d] <= 8'hf0;
		memory[16'h550e] <= 8'hb5;
		memory[16'h550f] <= 8'h3b;
		memory[16'h5510] <= 8'hcb;
		memory[16'h5511] <= 8'hef;
		memory[16'h5512] <= 8'hfd;
		memory[16'h5513] <= 8'h9b;
		memory[16'h5514] <= 8'hd1;
		memory[16'h5515] <= 8'hcd;
		memory[16'h5516] <= 8'h1f;
		memory[16'h5517] <= 8'hec;
		memory[16'h5518] <= 8'he3;
		memory[16'h5519] <= 8'hb9;
		memory[16'h551a] <= 8'h9e;
		memory[16'h551b] <= 8'h8e;
		memory[16'h551c] <= 8'h16;
		memory[16'h551d] <= 8'hc4;
		memory[16'h551e] <= 8'hd8;
		memory[16'h551f] <= 8'hbc;
		memory[16'h5520] <= 8'h99;
		memory[16'h5521] <= 8'h7f;
		memory[16'h5522] <= 8'h53;
		memory[16'h5523] <= 8'h14;
		memory[16'h5524] <= 8'hba;
		memory[16'h5525] <= 8'hd6;
		memory[16'h5526] <= 8'h26;
		memory[16'h5527] <= 8'h47;
		memory[16'h5528] <= 8'h2e;
		memory[16'h5529] <= 8'hbe;
		memory[16'h552a] <= 8'h37;
		memory[16'h552b] <= 8'h87;
		memory[16'h552c] <= 8'hae;
		memory[16'h552d] <= 8'hec;
		memory[16'h552e] <= 8'hc2;
		memory[16'h552f] <= 8'h79;
		memory[16'h5530] <= 8'hdb;
		memory[16'h5531] <= 8'hbf;
		memory[16'h5532] <= 8'h14;
		memory[16'h5533] <= 8'hac;
		memory[16'h5534] <= 8'h8d;
		memory[16'h5535] <= 8'h34;
		memory[16'h5536] <= 8'h98;
		memory[16'h5537] <= 8'h70;
		memory[16'h5538] <= 8'hed;
		memory[16'h5539] <= 8'h37;
		memory[16'h553a] <= 8'hfe;
		memory[16'h553b] <= 8'h3;
		memory[16'h553c] <= 8'hfb;
		memory[16'h553d] <= 8'hd6;
		memory[16'h553e] <= 8'hbf;
		memory[16'h553f] <= 8'h94;
		memory[16'h5540] <= 8'h55;
		memory[16'h5541] <= 8'h12;
		memory[16'h5542] <= 8'ha8;
		memory[16'h5543] <= 8'hf;
		memory[16'h5544] <= 8'he8;
		memory[16'h5545] <= 8'hce;
		memory[16'h5546] <= 8'h56;
		memory[16'h5547] <= 8'h17;
		memory[16'h5548] <= 8'h8d;
		memory[16'h5549] <= 8'h8d;
		memory[16'h554a] <= 8'h9e;
		memory[16'h554b] <= 8'h3b;
		memory[16'h554c] <= 8'h79;
		memory[16'h554d] <= 8'h60;
		memory[16'h554e] <= 8'hb5;
		memory[16'h554f] <= 8'h54;
		memory[16'h5550] <= 8'h1f;
		memory[16'h5551] <= 8'hc9;
		memory[16'h5552] <= 8'h0;
		memory[16'h5553] <= 8'hac;
		memory[16'h5554] <= 8'hfd;
		memory[16'h5555] <= 8'h99;
		memory[16'h5556] <= 8'h1c;
		memory[16'h5557] <= 8'hea;
		memory[16'h5558] <= 8'hd0;
		memory[16'h5559] <= 8'h1a;
		memory[16'h555a] <= 8'hee;
		memory[16'h555b] <= 8'hcb;
		memory[16'h555c] <= 8'hf0;
		memory[16'h555d] <= 8'had;
		memory[16'h555e] <= 8'h5f;
		memory[16'h555f] <= 8'h45;
		memory[16'h5560] <= 8'hc0;
		memory[16'h5561] <= 8'h7;
		memory[16'h5562] <= 8'h54;
		memory[16'h5563] <= 8'ha8;
		memory[16'h5564] <= 8'hd5;
		memory[16'h5565] <= 8'haa;
		memory[16'h5566] <= 8'hbf;
		memory[16'h5567] <= 8'h62;
		memory[16'h5568] <= 8'h37;
		memory[16'h5569] <= 8'h5d;
		memory[16'h556a] <= 8'h9e;
		memory[16'h556b] <= 8'hb0;
		memory[16'h556c] <= 8'hbd;
		memory[16'h556d] <= 8'h53;
		memory[16'h556e] <= 8'h4;
		memory[16'h556f] <= 8'hdd;
		memory[16'h5570] <= 8'h1c;
		memory[16'h5571] <= 8'h5;
		memory[16'h5572] <= 8'h89;
		memory[16'h5573] <= 8'h1a;
		memory[16'h5574] <= 8'h9e;
		memory[16'h5575] <= 8'ha6;
		memory[16'h5576] <= 8'h4;
		memory[16'h5577] <= 8'h6e;
		memory[16'h5578] <= 8'hc0;
		memory[16'h5579] <= 8'hf2;
		memory[16'h557a] <= 8'h39;
		memory[16'h557b] <= 8'hb1;
		memory[16'h557c] <= 8'ha0;
		memory[16'h557d] <= 8'h98;
		memory[16'h557e] <= 8'hf6;
		memory[16'h557f] <= 8'h60;
		memory[16'h5580] <= 8'h9f;
		memory[16'h5581] <= 8'h4b;
		memory[16'h5582] <= 8'h8;
		memory[16'h5583] <= 8'h74;
		memory[16'h5584] <= 8'hf5;
		memory[16'h5585] <= 8'hc8;
		memory[16'h5586] <= 8'hd7;
		memory[16'h5587] <= 8'h2d;
		memory[16'h5588] <= 8'h25;
		memory[16'h5589] <= 8'h75;
		memory[16'h558a] <= 8'hdd;
		memory[16'h558b] <= 8'he3;
		memory[16'h558c] <= 8'hc8;
		memory[16'h558d] <= 8'he2;
		memory[16'h558e] <= 8'hc0;
		memory[16'h558f] <= 8'he4;
		memory[16'h5590] <= 8'he7;
		memory[16'h5591] <= 8'h49;
		memory[16'h5592] <= 8'hfe;
		memory[16'h5593] <= 8'h85;
		memory[16'h5594] <= 8'hef;
		memory[16'h5595] <= 8'h3;
		memory[16'h5596] <= 8'hf3;
		memory[16'h5597] <= 8'hb0;
		memory[16'h5598] <= 8'hf5;
		memory[16'h5599] <= 8'h2c;
		memory[16'h559a] <= 8'h61;
		memory[16'h559b] <= 8'h95;
		memory[16'h559c] <= 8'hc4;
		memory[16'h559d] <= 8'h57;
		memory[16'h559e] <= 8'hf5;
		memory[16'h559f] <= 8'h63;
		memory[16'h55a0] <= 8'ha2;
		memory[16'h55a1] <= 8'hfe;
		memory[16'h55a2] <= 8'hd7;
		memory[16'h55a3] <= 8'h98;
		memory[16'h55a4] <= 8'hc6;
		memory[16'h55a5] <= 8'hae;
		memory[16'h55a6] <= 8'hc5;
		memory[16'h55a7] <= 8'heb;
		memory[16'h55a8] <= 8'h23;
		memory[16'h55a9] <= 8'ha2;
		memory[16'h55aa] <= 8'hce;
		memory[16'h55ab] <= 8'heb;
		memory[16'h55ac] <= 8'h84;
		memory[16'h55ad] <= 8'h8e;
		memory[16'h55ae] <= 8'hd0;
		memory[16'h55af] <= 8'h6b;
		memory[16'h55b0] <= 8'hd8;
		memory[16'h55b1] <= 8'hce;
		memory[16'h55b2] <= 8'hf0;
		memory[16'h55b3] <= 8'hc7;
		memory[16'h55b4] <= 8'hd1;
		memory[16'h55b5] <= 8'he3;
		memory[16'h55b6] <= 8'h77;
		memory[16'h55b7] <= 8'hc7;
		memory[16'h55b8] <= 8'hf;
		memory[16'h55b9] <= 8'hd8;
		memory[16'h55ba] <= 8'h5c;
		memory[16'h55bb] <= 8'hd3;
		memory[16'h55bc] <= 8'h30;
		memory[16'h55bd] <= 8'h52;
		memory[16'h55be] <= 8'h36;
		memory[16'h55bf] <= 8'hd2;
		memory[16'h55c0] <= 8'h50;
		memory[16'h55c1] <= 8'he;
		memory[16'h55c2] <= 8'h6a;
		memory[16'h55c3] <= 8'h16;
		memory[16'h55c4] <= 8'hbc;
		memory[16'h55c5] <= 8'h2f;
		memory[16'h55c6] <= 8'h1;
		memory[16'h55c7] <= 8'he0;
		memory[16'h55c8] <= 8'hd2;
		memory[16'h55c9] <= 8'hd0;
		memory[16'h55ca] <= 8'hcb;
		memory[16'h55cb] <= 8'h56;
		memory[16'h55cc] <= 8'h5e;
		memory[16'h55cd] <= 8'h9b;
		memory[16'h55ce] <= 8'hc2;
		memory[16'h55cf] <= 8'h36;
		memory[16'h55d0] <= 8'h6a;
		memory[16'h55d1] <= 8'hb2;
		memory[16'h55d2] <= 8'hfe;
		memory[16'h55d3] <= 8'h3b;
		memory[16'h55d4] <= 8'h96;
		memory[16'h55d5] <= 8'h75;
		memory[16'h55d6] <= 8'h2;
		memory[16'h55d7] <= 8'ha5;
		memory[16'h55d8] <= 8'h4e;
		memory[16'h55d9] <= 8'h5f;
		memory[16'h55da] <= 8'h79;
		memory[16'h55db] <= 8'h7e;
		memory[16'h55dc] <= 8'hb1;
		memory[16'h55dd] <= 8'haf;
		memory[16'h55de] <= 8'h50;
		memory[16'h55df] <= 8'h1;
		memory[16'h55e0] <= 8'hbd;
		memory[16'h55e1] <= 8'hbb;
		memory[16'h55e2] <= 8'h17;
		memory[16'h55e3] <= 8'h7a;
		memory[16'h55e4] <= 8'hea;
		memory[16'h55e5] <= 8'h18;
		memory[16'h55e6] <= 8'h5a;
		memory[16'h55e7] <= 8'hbc;
		memory[16'h55e8] <= 8'he8;
		memory[16'h55e9] <= 8'h25;
		memory[16'h55ea] <= 8'h13;
		memory[16'h55eb] <= 8'h47;
		memory[16'h55ec] <= 8'hc1;
		memory[16'h55ed] <= 8'hd5;
		memory[16'h55ee] <= 8'h7d;
		memory[16'h55ef] <= 8'h2b;
		memory[16'h55f0] <= 8'h87;
		memory[16'h55f1] <= 8'h7b;
		memory[16'h55f2] <= 8'h66;
		memory[16'h55f3] <= 8'h1d;
		memory[16'h55f4] <= 8'hf1;
		memory[16'h55f5] <= 8'h69;
		memory[16'h55f6] <= 8'hc3;
		memory[16'h55f7] <= 8'h3f;
		memory[16'h55f8] <= 8'hc8;
		memory[16'h55f9] <= 8'h3c;
		memory[16'h55fa] <= 8'hbd;
		memory[16'h55fb] <= 8'h79;
		memory[16'h55fc] <= 8'heb;
		memory[16'h55fd] <= 8'hd;
		memory[16'h55fe] <= 8'h7a;
		memory[16'h55ff] <= 8'ha9;
		memory[16'h5600] <= 8'hc8;
		memory[16'h5601] <= 8'h91;
		memory[16'h5602] <= 8'h23;
		memory[16'h5603] <= 8'hb3;
		memory[16'h5604] <= 8'ha9;
		memory[16'h5605] <= 8'h7d;
		memory[16'h5606] <= 8'h6f;
		memory[16'h5607] <= 8'h92;
		memory[16'h5608] <= 8'ha2;
		memory[16'h5609] <= 8'h82;
		memory[16'h560a] <= 8'hd9;
		memory[16'h560b] <= 8'h63;
		memory[16'h560c] <= 8'h57;
		memory[16'h560d] <= 8'h56;
		memory[16'h560e] <= 8'h8e;
		memory[16'h560f] <= 8'hdf;
		memory[16'h5610] <= 8'hd2;
		memory[16'h5611] <= 8'hf5;
		memory[16'h5612] <= 8'hfc;
		memory[16'h5613] <= 8'hc3;
		memory[16'h5614] <= 8'h5e;
		memory[16'h5615] <= 8'hbf;
		memory[16'h5616] <= 8'h2;
		memory[16'h5617] <= 8'h26;
		memory[16'h5618] <= 8'hfb;
		memory[16'h5619] <= 8'hbf;
		memory[16'h561a] <= 8'h9f;
		memory[16'h561b] <= 8'he7;
		memory[16'h561c] <= 8'hcc;
		memory[16'h561d] <= 8'h19;
		memory[16'h561e] <= 8'h90;
		memory[16'h561f] <= 8'h95;
		memory[16'h5620] <= 8'haa;
		memory[16'h5621] <= 8'hb3;
		memory[16'h5622] <= 8'h48;
		memory[16'h5623] <= 8'h53;
		memory[16'h5624] <= 8'h30;
		memory[16'h5625] <= 8'hb7;
		memory[16'h5626] <= 8'he5;
		memory[16'h5627] <= 8'hd2;
		memory[16'h5628] <= 8'h3a;
		memory[16'h5629] <= 8'hbe;
		memory[16'h562a] <= 8'h36;
		memory[16'h562b] <= 8'h91;
		memory[16'h562c] <= 8'h15;
		memory[16'h562d] <= 8'hc4;
		memory[16'h562e] <= 8'h70;
		memory[16'h562f] <= 8'he7;
		memory[16'h5630] <= 8'hb9;
		memory[16'h5631] <= 8'h6d;
		memory[16'h5632] <= 8'haa;
		memory[16'h5633] <= 8'h17;
		memory[16'h5634] <= 8'h2c;
		memory[16'h5635] <= 8'hac;
		memory[16'h5636] <= 8'h3d;
		memory[16'h5637] <= 8'h28;
		memory[16'h5638] <= 8'h6b;
		memory[16'h5639] <= 8'hdc;
		memory[16'h563a] <= 8'hf;
		memory[16'h563b] <= 8'h37;
		memory[16'h563c] <= 8'hf5;
		memory[16'h563d] <= 8'h9f;
		memory[16'h563e] <= 8'hcc;
		memory[16'h563f] <= 8'h9f;
		memory[16'h5640] <= 8'h52;
		memory[16'h5641] <= 8'h14;
		memory[16'h5642] <= 8'hf3;
		memory[16'h5643] <= 8'h82;
		memory[16'h5644] <= 8'hcc;
		memory[16'h5645] <= 8'hd8;
		memory[16'h5646] <= 8'h54;
		memory[16'h5647] <= 8'h6;
		memory[16'h5648] <= 8'h97;
		memory[16'h5649] <= 8'h8a;
		memory[16'h564a] <= 8'h97;
		memory[16'h564b] <= 8'hac;
		memory[16'h564c] <= 8'h4f;
		memory[16'h564d] <= 8'h8;
		memory[16'h564e] <= 8'h93;
		memory[16'h564f] <= 8'h8;
		memory[16'h5650] <= 8'h75;
		memory[16'h5651] <= 8'h3d;
		memory[16'h5652] <= 8'h20;
		memory[16'h5653] <= 8'ha1;
		memory[16'h5654] <= 8'he9;
		memory[16'h5655] <= 8'h5d;
		memory[16'h5656] <= 8'hc9;
		memory[16'h5657] <= 8'h54;
		memory[16'h5658] <= 8'h3a;
		memory[16'h5659] <= 8'hd8;
		memory[16'h565a] <= 8'h8b;
		memory[16'h565b] <= 8'h2f;
		memory[16'h565c] <= 8'h77;
		memory[16'h565d] <= 8'h58;
		memory[16'h565e] <= 8'hcf;
		memory[16'h565f] <= 8'hc9;
		memory[16'h5660] <= 8'h6c;
		memory[16'h5661] <= 8'hc2;
		memory[16'h5662] <= 8'h4b;
		memory[16'h5663] <= 8'h38;
		memory[16'h5664] <= 8'h9a;
		memory[16'h5665] <= 8'ha0;
		memory[16'h5666] <= 8'h3e;
		memory[16'h5667] <= 8'h31;
		memory[16'h5668] <= 8'h2a;
		memory[16'h5669] <= 8'hd6;
		memory[16'h566a] <= 8'hdd;
		memory[16'h566b] <= 8'h79;
		memory[16'h566c] <= 8'hde;
		memory[16'h566d] <= 8'h70;
		memory[16'h566e] <= 8'h82;
		memory[16'h566f] <= 8'h53;
		memory[16'h5670] <= 8'had;
		memory[16'h5671] <= 8'ha2;
		memory[16'h5672] <= 8'hf4;
		memory[16'h5673] <= 8'h96;
		memory[16'h5674] <= 8'hff;
		memory[16'h5675] <= 8'hbe;
		memory[16'h5676] <= 8'hea;
		memory[16'h5677] <= 8'h39;
		memory[16'h5678] <= 8'h96;
		memory[16'h5679] <= 8'h76;
		memory[16'h567a] <= 8'h69;
		memory[16'h567b] <= 8'he;
		memory[16'h567c] <= 8'hce;
		memory[16'h567d] <= 8'h38;
		memory[16'h567e] <= 8'hd7;
		memory[16'h567f] <= 8'h3a;
		memory[16'h5680] <= 8'hfa;
		memory[16'h5681] <= 8'h23;
		memory[16'h5682] <= 8'h73;
		memory[16'h5683] <= 8'h94;
		memory[16'h5684] <= 8'hc3;
		memory[16'h5685] <= 8'hb1;
		memory[16'h5686] <= 8'hc6;
		memory[16'h5687] <= 8'hed;
		memory[16'h5688] <= 8'h87;
		memory[16'h5689] <= 8'ha3;
		memory[16'h568a] <= 8'h67;
		memory[16'h568b] <= 8'h65;
		memory[16'h568c] <= 8'h14;
		memory[16'h568d] <= 8'he9;
		memory[16'h568e] <= 8'hb8;
		memory[16'h568f] <= 8'hc1;
		memory[16'h5690] <= 8'h8b;
		memory[16'h5691] <= 8'had;
		memory[16'h5692] <= 8'h58;
		memory[16'h5693] <= 8'h8a;
		memory[16'h5694] <= 8'h6b;
		memory[16'h5695] <= 8'h42;
		memory[16'h5696] <= 8'hc4;
		memory[16'h5697] <= 8'h1;
		memory[16'h5698] <= 8'hb8;
		memory[16'h5699] <= 8'h2d;
		memory[16'h569a] <= 8'hf;
		memory[16'h569b] <= 8'h86;
		memory[16'h569c] <= 8'h65;
		memory[16'h569d] <= 8'he7;
		memory[16'h569e] <= 8'hc1;
		memory[16'h569f] <= 8'h5f;
		memory[16'h56a0] <= 8'ha;
		memory[16'h56a1] <= 8'h34;
		memory[16'h56a2] <= 8'hf3;
		memory[16'h56a3] <= 8'hcd;
		memory[16'h56a4] <= 8'he5;
		memory[16'h56a5] <= 8'hb9;
		memory[16'h56a6] <= 8'hba;
		memory[16'h56a7] <= 8'h6d;
		memory[16'h56a8] <= 8'h5d;
		memory[16'h56a9] <= 8'h21;
		memory[16'h56aa] <= 8'hd2;
		memory[16'h56ab] <= 8'h71;
		memory[16'h56ac] <= 8'ha;
		memory[16'h56ad] <= 8'h8b;
		memory[16'h56ae] <= 8'h32;
		memory[16'h56af] <= 8'h95;
		memory[16'h56b0] <= 8'h38;
		memory[16'h56b1] <= 8'h8a;
		memory[16'h56b2] <= 8'h20;
		memory[16'h56b3] <= 8'ha3;
		memory[16'h56b4] <= 8'hcd;
		memory[16'h56b5] <= 8'he4;
		memory[16'h56b6] <= 8'ha4;
		memory[16'h56b7] <= 8'h85;
		memory[16'h56b8] <= 8'h11;
		memory[16'h56b9] <= 8'hb4;
		memory[16'h56ba] <= 8'hc;
		memory[16'h56bb] <= 8'h76;
		memory[16'h56bc] <= 8'h9b;
		memory[16'h56bd] <= 8'hcd;
		memory[16'h56be] <= 8'hd5;
		memory[16'h56bf] <= 8'ha5;
		memory[16'h56c0] <= 8'h1;
		memory[16'h56c1] <= 8'hc8;
		memory[16'h56c2] <= 8'h72;
		memory[16'h56c3] <= 8'he6;
		memory[16'h56c4] <= 8'h82;
		memory[16'h56c5] <= 8'h2c;
		memory[16'h56c6] <= 8'h53;
		memory[16'h56c7] <= 8'hdf;
		memory[16'h56c8] <= 8'h4e;
		memory[16'h56c9] <= 8'h26;
		memory[16'h56ca] <= 8'h50;
		memory[16'h56cb] <= 8'h58;
		memory[16'h56cc] <= 8'hb1;
		memory[16'h56cd] <= 8'h82;
		memory[16'h56ce] <= 8'hee;
		memory[16'h56cf] <= 8'he9;
		memory[16'h56d0] <= 8'hd;
		memory[16'h56d1] <= 8'he;
		memory[16'h56d2] <= 8'h8c;
		memory[16'h56d3] <= 8'hda;
		memory[16'h56d4] <= 8'hf2;
		memory[16'h56d5] <= 8'h30;
		memory[16'h56d6] <= 8'h5f;
		memory[16'h56d7] <= 8'h3;
		memory[16'h56d8] <= 8'he4;
		memory[16'h56d9] <= 8'h6b;
		memory[16'h56da] <= 8'h79;
		memory[16'h56db] <= 8'h7f;
		memory[16'h56dc] <= 8'h38;
		memory[16'h56dd] <= 8'h4e;
		memory[16'h56de] <= 8'h24;
		memory[16'h56df] <= 8'h39;
		memory[16'h56e0] <= 8'h16;
		memory[16'h56e1] <= 8'h96;
		memory[16'h56e2] <= 8'h20;
		memory[16'h56e3] <= 8'h98;
		memory[16'h56e4] <= 8'hc3;
		memory[16'h56e5] <= 8'h73;
		memory[16'h56e6] <= 8'h77;
		memory[16'h56e7] <= 8'h11;
		memory[16'h56e8] <= 8'h99;
		memory[16'h56e9] <= 8'hc7;
		memory[16'h56ea] <= 8'h69;
		memory[16'h56eb] <= 8'h4a;
		memory[16'h56ec] <= 8'h4a;
		memory[16'h56ed] <= 8'h57;
		memory[16'h56ee] <= 8'h33;
		memory[16'h56ef] <= 8'h57;
		memory[16'h56f0] <= 8'h65;
		memory[16'h56f1] <= 8'hbf;
		memory[16'h56f2] <= 8'h31;
		memory[16'h56f3] <= 8'h57;
		memory[16'h56f4] <= 8'hf0;
		memory[16'h56f5] <= 8'h90;
		memory[16'h56f6] <= 8'h5a;
		memory[16'h56f7] <= 8'hd4;
		memory[16'h56f8] <= 8'hfc;
		memory[16'h56f9] <= 8'hd3;
		memory[16'h56fa] <= 8'h54;
		memory[16'h56fb] <= 8'h34;
		memory[16'h56fc] <= 8'h21;
		memory[16'h56fd] <= 8'h78;
		memory[16'h56fe] <= 8'h6e;
		memory[16'h56ff] <= 8'h38;
		memory[16'h5700] <= 8'hf;
		memory[16'h5701] <= 8'h8e;
		memory[16'h5702] <= 8'hd0;
		memory[16'h5703] <= 8'hd2;
		memory[16'h5704] <= 8'h1;
		memory[16'h5705] <= 8'h48;
		memory[16'h5706] <= 8'he3;
		memory[16'h5707] <= 8'h9b;
		memory[16'h5708] <= 8'hf;
		memory[16'h5709] <= 8'h4c;
		memory[16'h570a] <= 8'he5;
		memory[16'h570b] <= 8'h59;
		memory[16'h570c] <= 8'ha4;
		memory[16'h570d] <= 8'h19;
		memory[16'h570e] <= 8'hb0;
		memory[16'h570f] <= 8'h9;
		memory[16'h5710] <= 8'hd8;
		memory[16'h5711] <= 8'he1;
		memory[16'h5712] <= 8'h61;
		memory[16'h5713] <= 8'hc8;
		memory[16'h5714] <= 8'h72;
		memory[16'h5715] <= 8'hbb;
		memory[16'h5716] <= 8'h9d;
		memory[16'h5717] <= 8'h6e;
		memory[16'h5718] <= 8'h8f;
		memory[16'h5719] <= 8'hf1;
		memory[16'h571a] <= 8'ha2;
		memory[16'h571b] <= 8'hb0;
		memory[16'h571c] <= 8'h69;
		memory[16'h571d] <= 8'h10;
		memory[16'h571e] <= 8'he8;
		memory[16'h571f] <= 8'h78;
		memory[16'h5720] <= 8'h9e;
		memory[16'h5721] <= 8'hb9;
		memory[16'h5722] <= 8'h4a;
		memory[16'h5723] <= 8'ha0;
		memory[16'h5724] <= 8'h1;
		memory[16'h5725] <= 8'h2d;
		memory[16'h5726] <= 8'h3b;
		memory[16'h5727] <= 8'h10;
		memory[16'h5728] <= 8'h7a;
		memory[16'h5729] <= 8'h20;
		memory[16'h572a] <= 8'h6a;
		memory[16'h572b] <= 8'h1e;
		memory[16'h572c] <= 8'h39;
		memory[16'h572d] <= 8'h1a;
		memory[16'h572e] <= 8'h27;
		memory[16'h572f] <= 8'h12;
		memory[16'h5730] <= 8'hfc;
		memory[16'h5731] <= 8'h88;
		memory[16'h5732] <= 8'hda;
		memory[16'h5733] <= 8'h6e;
		memory[16'h5734] <= 8'h44;
		memory[16'h5735] <= 8'h77;
		memory[16'h5736] <= 8'hdc;
		memory[16'h5737] <= 8'hd3;
		memory[16'h5738] <= 8'h68;
		memory[16'h5739] <= 8'h7e;
		memory[16'h573a] <= 8'h83;
		memory[16'h573b] <= 8'hd2;
		memory[16'h573c] <= 8'h8f;
		memory[16'h573d] <= 8'h6c;
		memory[16'h573e] <= 8'h4a;
		memory[16'h573f] <= 8'h2d;
		memory[16'h5740] <= 8'h25;
		memory[16'h5741] <= 8'h95;
		memory[16'h5742] <= 8'hcd;
		memory[16'h5743] <= 8'h26;
		memory[16'h5744] <= 8'hc2;
		memory[16'h5745] <= 8'h8;
		memory[16'h5746] <= 8'h36;
		memory[16'h5747] <= 8'h3c;
		memory[16'h5748] <= 8'h29;
		memory[16'h5749] <= 8'ha0;
		memory[16'h574a] <= 8'h5a;
		memory[16'h574b] <= 8'h62;
		memory[16'h574c] <= 8'hbb;
		memory[16'h574d] <= 8'h82;
		memory[16'h574e] <= 8'h74;
		memory[16'h574f] <= 8'hb7;
		memory[16'h5750] <= 8'ha;
		memory[16'h5751] <= 8'h4f;
		memory[16'h5752] <= 8'h25;
		memory[16'h5753] <= 8'h4e;
		memory[16'h5754] <= 8'hc6;
		memory[16'h5755] <= 8'h1;
		memory[16'h5756] <= 8'h21;
		memory[16'h5757] <= 8'h2f;
		memory[16'h5758] <= 8'h7f;
		memory[16'h5759] <= 8'ha5;
		memory[16'h575a] <= 8'h1;
		memory[16'h575b] <= 8'he;
		memory[16'h575c] <= 8'h11;
		memory[16'h575d] <= 8'h4b;
		memory[16'h575e] <= 8'h3c;
		memory[16'h575f] <= 8'h36;
		memory[16'h5760] <= 8'he0;
		memory[16'h5761] <= 8'h9;
		memory[16'h5762] <= 8'h5c;
		memory[16'h5763] <= 8'ha3;
		memory[16'h5764] <= 8'h12;
		memory[16'h5765] <= 8'h92;
		memory[16'h5766] <= 8'hdf;
		memory[16'h5767] <= 8'h3b;
		memory[16'h5768] <= 8'h33;
		memory[16'h5769] <= 8'h3a;
		memory[16'h576a] <= 8'h9d;
		memory[16'h576b] <= 8'hee;
		memory[16'h576c] <= 8'hbc;
		memory[16'h576d] <= 8'h12;
		memory[16'h576e] <= 8'ha5;
		memory[16'h576f] <= 8'hc6;
		memory[16'h5770] <= 8'h61;
		memory[16'h5771] <= 8'hca;
		memory[16'h5772] <= 8'h15;
		memory[16'h5773] <= 8'h27;
		memory[16'h5774] <= 8'hcb;
		memory[16'h5775] <= 8'h36;
		memory[16'h5776] <= 8'h56;
		memory[16'h5777] <= 8'h4a;
		memory[16'h5778] <= 8'hdb;
		memory[16'h5779] <= 8'h57;
		memory[16'h577a] <= 8'h59;
		memory[16'h577b] <= 8'hec;
		memory[16'h577c] <= 8'ha3;
		memory[16'h577d] <= 8'h95;
		memory[16'h577e] <= 8'h22;
		memory[16'h577f] <= 8'h83;
		memory[16'h5780] <= 8'h9e;
		memory[16'h5781] <= 8'h7e;
		memory[16'h5782] <= 8'h26;
		memory[16'h5783] <= 8'hb0;
		memory[16'h5784] <= 8'h11;
		memory[16'h5785] <= 8'h6;
		memory[16'h5786] <= 8'heb;
		memory[16'h5787] <= 8'h44;
		memory[16'h5788] <= 8'h40;
		memory[16'h5789] <= 8'h89;
		memory[16'h578a] <= 8'h32;
		memory[16'h578b] <= 8'hfc;
		memory[16'h578c] <= 8'h9b;
		memory[16'h578d] <= 8'hd7;
		memory[16'h578e] <= 8'hc2;
		memory[16'h578f] <= 8'hfc;
		memory[16'h5790] <= 8'ha1;
		memory[16'h5791] <= 8'hd7;
		memory[16'h5792] <= 8'h23;
		memory[16'h5793] <= 8'h6c;
		memory[16'h5794] <= 8'he;
		memory[16'h5795] <= 8'h7a;
		memory[16'h5796] <= 8'hb6;
		memory[16'h5797] <= 8'he9;
		memory[16'h5798] <= 8'hd1;
		memory[16'h5799] <= 8'hf;
		memory[16'h579a] <= 8'hd6;
		memory[16'h579b] <= 8'h74;
		memory[16'h579c] <= 8'ha4;
		memory[16'h579d] <= 8'hf8;
		memory[16'h579e] <= 8'hf8;
		memory[16'h579f] <= 8'h43;
		memory[16'h57a0] <= 8'h77;
		memory[16'h57a1] <= 8'h1e;
		memory[16'h57a2] <= 8'hf3;
		memory[16'h57a3] <= 8'h88;
		memory[16'h57a4] <= 8'h24;
		memory[16'h57a5] <= 8'hdf;
		memory[16'h57a6] <= 8'hcc;
		memory[16'h57a7] <= 8'h64;
		memory[16'h57a8] <= 8'h68;
		memory[16'h57a9] <= 8'hfe;
		memory[16'h57aa] <= 8'h60;
		memory[16'h57ab] <= 8'h3;
		memory[16'h57ac] <= 8'hd5;
		memory[16'h57ad] <= 8'h23;
		memory[16'h57ae] <= 8'hff;
		memory[16'h57af] <= 8'h76;
		memory[16'h57b0] <= 8'hfa;
		memory[16'h57b1] <= 8'h22;
		memory[16'h57b2] <= 8'he2;
		memory[16'h57b3] <= 8'h8;
		memory[16'h57b4] <= 8'h9c;
		memory[16'h57b5] <= 8'h98;
		memory[16'h57b6] <= 8'hf2;
		memory[16'h57b7] <= 8'h6e;
		memory[16'h57b8] <= 8'ha8;
		memory[16'h57b9] <= 8'hc8;
		memory[16'h57ba] <= 8'he2;
		memory[16'h57bb] <= 8'h4c;
		memory[16'h57bc] <= 8'hc0;
		memory[16'h57bd] <= 8'hda;
		memory[16'h57be] <= 8'h8f;
		memory[16'h57bf] <= 8'h37;
		memory[16'h57c0] <= 8'hf9;
		memory[16'h57c1] <= 8'h83;
		memory[16'h57c2] <= 8'hbf;
		memory[16'h57c3] <= 8'h1d;
		memory[16'h57c4] <= 8'h62;
		memory[16'h57c5] <= 8'h8b;
		memory[16'h57c6] <= 8'h82;
		memory[16'h57c7] <= 8'hca;
		memory[16'h57c8] <= 8'h89;
		memory[16'h57c9] <= 8'he2;
		memory[16'h57ca] <= 8'hcd;
		memory[16'h57cb] <= 8'h5e;
		memory[16'h57cc] <= 8'h5;
		memory[16'h57cd] <= 8'hcc;
		memory[16'h57ce] <= 8'hd4;
		memory[16'h57cf] <= 8'h0;
		memory[16'h57d0] <= 8'hee;
		memory[16'h57d1] <= 8'hb6;
		memory[16'h57d2] <= 8'h8;
		memory[16'h57d3] <= 8'h8b;
		memory[16'h57d4] <= 8'h4f;
		memory[16'h57d5] <= 8'hfa;
		memory[16'h57d6] <= 8'hf9;
		memory[16'h57d7] <= 8'hf7;
		memory[16'h57d8] <= 8'hc2;
		memory[16'h57d9] <= 8'hdb;
		memory[16'h57da] <= 8'h43;
		memory[16'h57db] <= 8'h83;
		memory[16'h57dc] <= 8'hb6;
		memory[16'h57dd] <= 8'hd3;
		memory[16'h57de] <= 8'hba;
		memory[16'h57df] <= 8'haf;
		memory[16'h57e0] <= 8'h56;
		memory[16'h57e1] <= 8'h7a;
		memory[16'h57e2] <= 8'hcc;
		memory[16'h57e3] <= 8'hb8;
		memory[16'h57e4] <= 8'h5;
		memory[16'h57e5] <= 8'h4e;
		memory[16'h57e6] <= 8'h82;
		memory[16'h57e7] <= 8'h8f;
		memory[16'h57e8] <= 8'h31;
		memory[16'h57e9] <= 8'h4f;
		memory[16'h57ea] <= 8'hed;
		memory[16'h57eb] <= 8'h36;
		memory[16'h57ec] <= 8'h1b;
		memory[16'h57ed] <= 8'hc2;
		memory[16'h57ee] <= 8'h36;
		memory[16'h57ef] <= 8'h9;
		memory[16'h57f0] <= 8'h78;
		memory[16'h57f1] <= 8'h3f;
		memory[16'h57f2] <= 8'h94;
		memory[16'h57f3] <= 8'hc7;
		memory[16'h57f4] <= 8'h39;
		memory[16'h57f5] <= 8'h8d;
		memory[16'h57f6] <= 8'hbe;
		memory[16'h57f7] <= 8'hfc;
		memory[16'h57f8] <= 8'h69;
		memory[16'h57f9] <= 8'h2;
		memory[16'h57fa] <= 8'h7f;
		memory[16'h57fb] <= 8'h1f;
		memory[16'h57fc] <= 8'hd5;
		memory[16'h57fd] <= 8'h39;
		memory[16'h57fe] <= 8'hce;
		memory[16'h57ff] <= 8'h2b;
		memory[16'h5800] <= 8'hb3;
		memory[16'h5801] <= 8'h9a;
		memory[16'h5802] <= 8'he3;
		memory[16'h5803] <= 8'hb9;
		memory[16'h5804] <= 8'he9;
		memory[16'h5805] <= 8'h65;
		memory[16'h5806] <= 8'h48;
		memory[16'h5807] <= 8'h1a;
		memory[16'h5808] <= 8'hb4;
		memory[16'h5809] <= 8'h35;
		memory[16'h580a] <= 8'h50;
		memory[16'h580b] <= 8'hcf;
		memory[16'h580c] <= 8'hf7;
		memory[16'h580d] <= 8'h87;
		memory[16'h580e] <= 8'hd8;
		memory[16'h580f] <= 8'h70;
		memory[16'h5810] <= 8'hc6;
		memory[16'h5811] <= 8'h6d;
		memory[16'h5812] <= 8'h37;
		memory[16'h5813] <= 8'hff;
		memory[16'h5814] <= 8'hfa;
		memory[16'h5815] <= 8'hf6;
		memory[16'h5816] <= 8'hfb;
		memory[16'h5817] <= 8'h63;
		memory[16'h5818] <= 8'hf8;
		memory[16'h5819] <= 8'h7a;
		memory[16'h581a] <= 8'h82;
		memory[16'h581b] <= 8'hcd;
		memory[16'h581c] <= 8'hb4;
		memory[16'h581d] <= 8'h50;
		memory[16'h581e] <= 8'hf8;
		memory[16'h581f] <= 8'h67;
		memory[16'h5820] <= 8'heb;
		memory[16'h5821] <= 8'hdb;
		memory[16'h5822] <= 8'h20;
		memory[16'h5823] <= 8'hd4;
		memory[16'h5824] <= 8'h40;
		memory[16'h5825] <= 8'h68;
		memory[16'h5826] <= 8'hee;
		memory[16'h5827] <= 8'hf4;
		memory[16'h5828] <= 8'h9e;
		memory[16'h5829] <= 8'h3e;
		memory[16'h582a] <= 8'hc3;
		memory[16'h582b] <= 8'h95;
		memory[16'h582c] <= 8'hc5;
		memory[16'h582d] <= 8'h9b;
		memory[16'h582e] <= 8'h5;
		memory[16'h582f] <= 8'h8b;
		memory[16'h5830] <= 8'h8;
		memory[16'h5831] <= 8'h3d;
		memory[16'h5832] <= 8'h8b;
		memory[16'h5833] <= 8'h3;
		memory[16'h5834] <= 8'h33;
		memory[16'h5835] <= 8'h86;
		memory[16'h5836] <= 8'h66;
		memory[16'h5837] <= 8'h2b;
		memory[16'h5838] <= 8'h1;
		memory[16'h5839] <= 8'he9;
		memory[16'h583a] <= 8'hf8;
		memory[16'h583b] <= 8'hb5;
		memory[16'h583c] <= 8'h39;
		memory[16'h583d] <= 8'hf0;
		memory[16'h583e] <= 8'h1c;
		memory[16'h583f] <= 8'h24;
		memory[16'h5840] <= 8'hcb;
		memory[16'h5841] <= 8'h3d;
		memory[16'h5842] <= 8'hf8;
		memory[16'h5843] <= 8'hb;
		memory[16'h5844] <= 8'ha5;
		memory[16'h5845] <= 8'he6;
		memory[16'h5846] <= 8'hff;
		memory[16'h5847] <= 8'h43;
		memory[16'h5848] <= 8'h25;
		memory[16'h5849] <= 8'hc2;
		memory[16'h584a] <= 8'hd9;
		memory[16'h584b] <= 8'hea;
		memory[16'h584c] <= 8'h5d;
		memory[16'h584d] <= 8'hde;
		memory[16'h584e] <= 8'h76;
		memory[16'h584f] <= 8'h66;
		memory[16'h5850] <= 8'h1b;
		memory[16'h5851] <= 8'h1;
		memory[16'h5852] <= 8'h69;
		memory[16'h5853] <= 8'h4e;
		memory[16'h5854] <= 8'h87;
		memory[16'h5855] <= 8'hcf;
		memory[16'h5856] <= 8'h79;
		memory[16'h5857] <= 8'h88;
		memory[16'h5858] <= 8'hb8;
		memory[16'h5859] <= 8'h71;
		memory[16'h585a] <= 8'h3d;
		memory[16'h585b] <= 8'hf2;
		memory[16'h585c] <= 8'h61;
		memory[16'h585d] <= 8'h5a;
		memory[16'h585e] <= 8'h16;
		memory[16'h585f] <= 8'h2c;
		memory[16'h5860] <= 8'h97;
		memory[16'h5861] <= 8'hf;
		memory[16'h5862] <= 8'h37;
		memory[16'h5863] <= 8'h3c;
		memory[16'h5864] <= 8'hf5;
		memory[16'h5865] <= 8'h36;
		memory[16'h5866] <= 8'h80;
		memory[16'h5867] <= 8'h1a;
		memory[16'h5868] <= 8'hf8;
		memory[16'h5869] <= 8'h59;
		memory[16'h586a] <= 8'h5;
		memory[16'h586b] <= 8'h56;
		memory[16'h586c] <= 8'h37;
		memory[16'h586d] <= 8'h7b;
		memory[16'h586e] <= 8'hbc;
		memory[16'h586f] <= 8'h53;
		memory[16'h5870] <= 8'h7c;
		memory[16'h5871] <= 8'h25;
		memory[16'h5872] <= 8'ha1;
		memory[16'h5873] <= 8'h3;
		memory[16'h5874] <= 8'hf4;
		memory[16'h5875] <= 8'h1b;
		memory[16'h5876] <= 8'h8c;
		memory[16'h5877] <= 8'had;
		memory[16'h5878] <= 8'h8c;
		memory[16'h5879] <= 8'hc9;
		memory[16'h587a] <= 8'h9f;
		memory[16'h587b] <= 8'hee;
		memory[16'h587c] <= 8'h23;
		memory[16'h587d] <= 8'hb5;
		memory[16'h587e] <= 8'h1a;
		memory[16'h587f] <= 8'hba;
		memory[16'h5880] <= 8'hc4;
		memory[16'h5881] <= 8'h52;
		memory[16'h5882] <= 8'hf7;
		memory[16'h5883] <= 8'hba;
		memory[16'h5884] <= 8'h88;
		memory[16'h5885] <= 8'h77;
		memory[16'h5886] <= 8'hd4;
		memory[16'h5887] <= 8'h81;
		memory[16'h5888] <= 8'hd0;
		memory[16'h5889] <= 8'hd9;
		memory[16'h588a] <= 8'hd7;
		memory[16'h588b] <= 8'h7;
		memory[16'h588c] <= 8'h54;
		memory[16'h588d] <= 8'h93;
		memory[16'h588e] <= 8'h5a;
		memory[16'h588f] <= 8'hd0;
		memory[16'h5890] <= 8'hb8;
		memory[16'h5891] <= 8'hfc;
		memory[16'h5892] <= 8'hd4;
		memory[16'h5893] <= 8'hac;
		memory[16'h5894] <= 8'h17;
		memory[16'h5895] <= 8'h60;
		memory[16'h5896] <= 8'h59;
		memory[16'h5897] <= 8'ha3;
		memory[16'h5898] <= 8'h29;
		memory[16'h5899] <= 8'hf8;
		memory[16'h589a] <= 8'h91;
		memory[16'h589b] <= 8'h4d;
		memory[16'h589c] <= 8'hae;
		memory[16'h589d] <= 8'hac;
		memory[16'h589e] <= 8'h7;
		memory[16'h589f] <= 8'h72;
		memory[16'h58a0] <= 8'hfe;
		memory[16'h58a1] <= 8'hfe;
		memory[16'h58a2] <= 8'h2c;
		memory[16'h58a3] <= 8'h86;
		memory[16'h58a4] <= 8'h75;
		memory[16'h58a5] <= 8'h1;
		memory[16'h58a6] <= 8'h7;
		memory[16'h58a7] <= 8'h45;
		memory[16'h58a8] <= 8'hda;
		memory[16'h58a9] <= 8'hde;
		memory[16'h58aa] <= 8'h4d;
		memory[16'h58ab] <= 8'h2f;
		memory[16'h58ac] <= 8'h71;
		memory[16'h58ad] <= 8'ha7;
		memory[16'h58ae] <= 8'hff;
		memory[16'h58af] <= 8'h29;
		memory[16'h58b0] <= 8'ha3;
		memory[16'h58b1] <= 8'hd3;
		memory[16'h58b2] <= 8'hd6;
		memory[16'h58b3] <= 8'hba;
		memory[16'h58b4] <= 8'h33;
		memory[16'h58b5] <= 8'h2f;
		memory[16'h58b6] <= 8'h5e;
		memory[16'h58b7] <= 8'h5d;
		memory[16'h58b8] <= 8'h28;
		memory[16'h58b9] <= 8'hef;
		memory[16'h58ba] <= 8'haa;
		memory[16'h58bb] <= 8'hd6;
		memory[16'h58bc] <= 8'h9b;
		memory[16'h58bd] <= 8'hb1;
		memory[16'h58be] <= 8'h48;
		memory[16'h58bf] <= 8'h99;
		memory[16'h58c0] <= 8'hb0;
		memory[16'h58c1] <= 8'h75;
		memory[16'h58c2] <= 8'h20;
		memory[16'h58c3] <= 8'h25;
		memory[16'h58c4] <= 8'h76;
		memory[16'h58c5] <= 8'h27;
		memory[16'h58c6] <= 8'h6b;
		memory[16'h58c7] <= 8'h50;
		memory[16'h58c8] <= 8'h6;
		memory[16'h58c9] <= 8'hb8;
		memory[16'h58ca] <= 8'h7f;
		memory[16'h58cb] <= 8'h77;
		memory[16'h58cc] <= 8'h5f;
		memory[16'h58cd] <= 8'h7f;
		memory[16'h58ce] <= 8'ha1;
		memory[16'h58cf] <= 8'h3;
		memory[16'h58d0] <= 8'h52;
		memory[16'h58d1] <= 8'h77;
		memory[16'h58d2] <= 8'hbd;
		memory[16'h58d3] <= 8'h86;
		memory[16'h58d4] <= 8'ha6;
		memory[16'h58d5] <= 8'h1b;
		memory[16'h58d6] <= 8'he3;
		memory[16'h58d7] <= 8'hce;
		memory[16'h58d8] <= 8'hb;
		memory[16'h58d9] <= 8'h8d;
		memory[16'h58da] <= 8'ha4;
		memory[16'h58db] <= 8'ha6;
		memory[16'h58dc] <= 8'h3e;
		memory[16'h58dd] <= 8'hed;
		memory[16'h58de] <= 8'h40;
		memory[16'h58df] <= 8'hee;
		memory[16'h58e0] <= 8'h62;
		memory[16'h58e1] <= 8'h60;
		memory[16'h58e2] <= 8'h14;
		memory[16'h58e3] <= 8'hd8;
		memory[16'h58e4] <= 8'h87;
		memory[16'h58e5] <= 8'h7f;
		memory[16'h58e6] <= 8'h28;
		memory[16'h58e7] <= 8'h8d;
		memory[16'h58e8] <= 8'h37;
		memory[16'h58e9] <= 8'ha8;
		memory[16'h58ea] <= 8'h5;
		memory[16'h58eb] <= 8'h96;
		memory[16'h58ec] <= 8'h27;
		memory[16'h58ed] <= 8'ha6;
		memory[16'h58ee] <= 8'h99;
		memory[16'h58ef] <= 8'h79;
		memory[16'h58f0] <= 8'h1d;
		memory[16'h58f1] <= 8'h57;
		memory[16'h58f2] <= 8'hff;
		memory[16'h58f3] <= 8'hc3;
		memory[16'h58f4] <= 8'h72;
		memory[16'h58f5] <= 8'he2;
		memory[16'h58f6] <= 8'h92;
		memory[16'h58f7] <= 8'h7d;
		memory[16'h58f8] <= 8'h6f;
		memory[16'h58f9] <= 8'h36;
		memory[16'h58fa] <= 8'h24;
		memory[16'h58fb] <= 8'hae;
		memory[16'h58fc] <= 8'h23;
		memory[16'h58fd] <= 8'h64;
		memory[16'h58fe] <= 8'h9c;
		memory[16'h58ff] <= 8'h85;
		memory[16'h5900] <= 8'hc4;
		memory[16'h5901] <= 8'hb0;
		memory[16'h5902] <= 8'h5d;
		memory[16'h5903] <= 8'h4b;
		memory[16'h5904] <= 8'h2f;
		memory[16'h5905] <= 8'h86;
		memory[16'h5906] <= 8'hd9;
		memory[16'h5907] <= 8'h66;
		memory[16'h5908] <= 8'h2e;
		memory[16'h5909] <= 8'hde;
		memory[16'h590a] <= 8'hfd;
		memory[16'h590b] <= 8'h55;
		memory[16'h590c] <= 8'h84;
		memory[16'h590d] <= 8'h96;
		memory[16'h590e] <= 8'hce;
		memory[16'h590f] <= 8'ha1;
		memory[16'h5910] <= 8'hed;
		memory[16'h5911] <= 8'hce;
		memory[16'h5912] <= 8'h64;
		memory[16'h5913] <= 8'h60;
		memory[16'h5914] <= 8'hb0;
		memory[16'h5915] <= 8'hf6;
		memory[16'h5916] <= 8'hdd;
		memory[16'h5917] <= 8'h20;
		memory[16'h5918] <= 8'h2d;
		memory[16'h5919] <= 8'h1;
		memory[16'h591a] <= 8'hce;
		memory[16'h591b] <= 8'h50;
		memory[16'h591c] <= 8'h65;
		memory[16'h591d] <= 8'h6a;
		memory[16'h591e] <= 8'hd6;
		memory[16'h591f] <= 8'h29;
		memory[16'h5920] <= 8'h1b;
		memory[16'h5921] <= 8'h33;
		memory[16'h5922] <= 8'h75;
		memory[16'h5923] <= 8'h4a;
		memory[16'h5924] <= 8'hb9;
		memory[16'h5925] <= 8'h4e;
		memory[16'h5926] <= 8'hb1;
		memory[16'h5927] <= 8'he7;
		memory[16'h5928] <= 8'h2c;
		memory[16'h5929] <= 8'hae;
		memory[16'h592a] <= 8'h3c;
		memory[16'h592b] <= 8'hb0;
		memory[16'h592c] <= 8'h44;
		memory[16'h592d] <= 8'hb;
		memory[16'h592e] <= 8'h51;
		memory[16'h592f] <= 8'h32;
		memory[16'h5930] <= 8'hd9;
		memory[16'h5931] <= 8'hb5;
		memory[16'h5932] <= 8'h92;
		memory[16'h5933] <= 8'h89;
		memory[16'h5934] <= 8'hac;
		memory[16'h5935] <= 8'h6f;
		memory[16'h5936] <= 8'ha9;
		memory[16'h5937] <= 8'hd9;
		memory[16'h5938] <= 8'h71;
		memory[16'h5939] <= 8'h77;
		memory[16'h593a] <= 8'h29;
		memory[16'h593b] <= 8'hd6;
		memory[16'h593c] <= 8'he2;
		memory[16'h593d] <= 8'hff;
		memory[16'h593e] <= 8'h0;
		memory[16'h593f] <= 8'hfd;
		memory[16'h5940] <= 8'h33;
		memory[16'h5941] <= 8'h75;
		memory[16'h5942] <= 8'h47;
		memory[16'h5943] <= 8'hec;
		memory[16'h5944] <= 8'hc3;
		memory[16'h5945] <= 8'hf8;
		memory[16'h5946] <= 8'hd4;
		memory[16'h5947] <= 8'hef;
		memory[16'h5948] <= 8'ha6;
		memory[16'h5949] <= 8'h10;
		memory[16'h594a] <= 8'h9f;
		memory[16'h594b] <= 8'heb;
		memory[16'h594c] <= 8'h1b;
		memory[16'h594d] <= 8'hf0;
		memory[16'h594e] <= 8'h1d;
		memory[16'h594f] <= 8'hf4;
		memory[16'h5950] <= 8'ha5;
		memory[16'h5951] <= 8'haf;
		memory[16'h5952] <= 8'h7e;
		memory[16'h5953] <= 8'h51;
		memory[16'h5954] <= 8'h1e;
		memory[16'h5955] <= 8'h27;
		memory[16'h5956] <= 8'h2a;
		memory[16'h5957] <= 8'h8f;
		memory[16'h5958] <= 8'h9f;
		memory[16'h5959] <= 8'h54;
		memory[16'h595a] <= 8'h66;
		memory[16'h595b] <= 8'h81;
		memory[16'h595c] <= 8'h53;
		memory[16'h595d] <= 8'h66;
		memory[16'h595e] <= 8'h7e;
		memory[16'h595f] <= 8'h86;
		memory[16'h5960] <= 8'hdb;
		memory[16'h5961] <= 8'hc5;
		memory[16'h5962] <= 8'h73;
		memory[16'h5963] <= 8'h9e;
		memory[16'h5964] <= 8'hbe;
		memory[16'h5965] <= 8'h47;
		memory[16'h5966] <= 8'h8d;
		memory[16'h5967] <= 8'h64;
		memory[16'h5968] <= 8'h57;
		memory[16'h5969] <= 8'h2c;
		memory[16'h596a] <= 8'h4f;
		memory[16'h596b] <= 8'h73;
		memory[16'h596c] <= 8'h1c;
		memory[16'h596d] <= 8'h6c;
		memory[16'h596e] <= 8'h67;
		memory[16'h596f] <= 8'hc1;
		memory[16'h5970] <= 8'h1b;
		memory[16'h5971] <= 8'he5;
		memory[16'h5972] <= 8'h13;
		memory[16'h5973] <= 8'h3a;
		memory[16'h5974] <= 8'hd;
		memory[16'h5975] <= 8'h3d;
		memory[16'h5976] <= 8'hc9;
		memory[16'h5977] <= 8'hac;
		memory[16'h5978] <= 8'h91;
		memory[16'h5979] <= 8'h2f;
		memory[16'h597a] <= 8'h2d;
		memory[16'h597b] <= 8'he5;
		memory[16'h597c] <= 8'h95;
		memory[16'h597d] <= 8'hab;
		memory[16'h597e] <= 8'h6b;
		memory[16'h597f] <= 8'h70;
		memory[16'h5980] <= 8'h70;
		memory[16'h5981] <= 8'hde;
		memory[16'h5982] <= 8'he;
		memory[16'h5983] <= 8'h2e;
		memory[16'h5984] <= 8'h25;
		memory[16'h5985] <= 8'h9b;
		memory[16'h5986] <= 8'h93;
		memory[16'h5987] <= 8'h7d;
		memory[16'h5988] <= 8'hc7;
		memory[16'h5989] <= 8'he2;
		memory[16'h598a] <= 8'hf0;
		memory[16'h598b] <= 8'he3;
		memory[16'h598c] <= 8'h4f;
		memory[16'h598d] <= 8'h57;
		memory[16'h598e] <= 8'ha5;
		memory[16'h598f] <= 8'h6a;
		memory[16'h5990] <= 8'h3d;
		memory[16'h5991] <= 8'hb8;
		memory[16'h5992] <= 8'ha4;
		memory[16'h5993] <= 8'h4a;
		memory[16'h5994] <= 8'hf5;
		memory[16'h5995] <= 8'h6e;
		memory[16'h5996] <= 8'hf6;
		memory[16'h5997] <= 8'h87;
		memory[16'h5998] <= 8'h9d;
		memory[16'h5999] <= 8'h23;
		memory[16'h599a] <= 8'h6c;
		memory[16'h599b] <= 8'h33;
		memory[16'h599c] <= 8'hce;
		memory[16'h599d] <= 8'hd7;
		memory[16'h599e] <= 8'ha3;
		memory[16'h599f] <= 8'h3e;
		memory[16'h59a0] <= 8'hb6;
		memory[16'h59a1] <= 8'hb2;
		memory[16'h59a2] <= 8'h6d;
		memory[16'h59a3] <= 8'hdb;
		memory[16'h59a4] <= 8'h4d;
		memory[16'h59a5] <= 8'h0;
		memory[16'h59a6] <= 8'h58;
		memory[16'h59a7] <= 8'h15;
		memory[16'h59a8] <= 8'he2;
		memory[16'h59a9] <= 8'h48;
		memory[16'h59aa] <= 8'hf8;
		memory[16'h59ab] <= 8'h31;
		memory[16'h59ac] <= 8'ha0;
		memory[16'h59ad] <= 8'h9d;
		memory[16'h59ae] <= 8'h9c;
		memory[16'h59af] <= 8'hdd;
		memory[16'h59b0] <= 8'h55;
		memory[16'h59b1] <= 8'h40;
		memory[16'h59b2] <= 8'h27;
		memory[16'h59b3] <= 8'h4b;
		memory[16'h59b4] <= 8'hae;
		memory[16'h59b5] <= 8'h1d;
		memory[16'h59b6] <= 8'hd2;
		memory[16'h59b7] <= 8'h4c;
		memory[16'h59b8] <= 8'h40;
		memory[16'h59b9] <= 8'h3e;
		memory[16'h59ba] <= 8'h7f;
		memory[16'h59bb] <= 8'he;
		memory[16'h59bc] <= 8'h15;
		memory[16'h59bd] <= 8'h22;
		memory[16'h59be] <= 8'h4c;
		memory[16'h59bf] <= 8'hcb;
		memory[16'h59c0] <= 8'hd4;
		memory[16'h59c1] <= 8'hb9;
		memory[16'h59c2] <= 8'ha7;
		memory[16'h59c3] <= 8'h22;
		memory[16'h59c4] <= 8'hb9;
		memory[16'h59c5] <= 8'hff;
		memory[16'h59c6] <= 8'h37;
		memory[16'h59c7] <= 8'h9c;
		memory[16'h59c8] <= 8'h48;
		memory[16'h59c9] <= 8'h2f;
		memory[16'h59ca] <= 8'hcd;
		memory[16'h59cb] <= 8'he8;
		memory[16'h59cc] <= 8'hcd;
		memory[16'h59cd] <= 8'h69;
		memory[16'h59ce] <= 8'hc5;
		memory[16'h59cf] <= 8'h22;
		memory[16'h59d0] <= 8'haa;
		memory[16'h59d1] <= 8'hec;
		memory[16'h59d2] <= 8'h6d;
		memory[16'h59d3] <= 8'h58;
		memory[16'h59d4] <= 8'h9;
		memory[16'h59d5] <= 8'h3f;
		memory[16'h59d6] <= 8'ha4;
		memory[16'h59d7] <= 8'h49;
		memory[16'h59d8] <= 8'h7d;
		memory[16'h59d9] <= 8'h23;
		memory[16'h59da] <= 8'h57;
		memory[16'h59db] <= 8'h93;
		memory[16'h59dc] <= 8'h46;
		memory[16'h59dd] <= 8'ha3;
		memory[16'h59de] <= 8'h5e;
		memory[16'h59df] <= 8'h1a;
		memory[16'h59e0] <= 8'h5d;
		memory[16'h59e1] <= 8'h5;
		memory[16'h59e2] <= 8'h3c;
		memory[16'h59e3] <= 8'h16;
		memory[16'h59e4] <= 8'h5;
		memory[16'h59e5] <= 8'h73;
		memory[16'h59e6] <= 8'hb2;
		memory[16'h59e7] <= 8'h4d;
		memory[16'h59e8] <= 8'ha3;
		memory[16'h59e9] <= 8'h80;
		memory[16'h59ea] <= 8'h35;
		memory[16'h59eb] <= 8'h70;
		memory[16'h59ec] <= 8'he9;
		memory[16'h59ed] <= 8'hfa;
		memory[16'h59ee] <= 8'h92;
		memory[16'h59ef] <= 8'h93;
		memory[16'h59f0] <= 8'he6;
		memory[16'h59f1] <= 8'h0;
		memory[16'h59f2] <= 8'hec;
		memory[16'h59f3] <= 8'hef;
		memory[16'h59f4] <= 8'h3f;
		memory[16'h59f5] <= 8'h90;
		memory[16'h59f6] <= 8'h38;
		memory[16'h59f7] <= 8'hbd;
		memory[16'h59f8] <= 8'hb4;
		memory[16'h59f9] <= 8'h8f;
		memory[16'h59fa] <= 8'h50;
		memory[16'h59fb] <= 8'hfa;
		memory[16'h59fc] <= 8'h32;
		memory[16'h59fd] <= 8'hae;
		memory[16'h59fe] <= 8'h14;
		memory[16'h59ff] <= 8'h8f;
		memory[16'h5a00] <= 8'hb4;
		memory[16'h5a01] <= 8'h51;
		memory[16'h5a02] <= 8'ha6;
		memory[16'h5a03] <= 8'hb9;
		memory[16'h5a04] <= 8'hc4;
		memory[16'h5a05] <= 8'h58;
		memory[16'h5a06] <= 8'h6;
		memory[16'h5a07] <= 8'h67;
		memory[16'h5a08] <= 8'hd8;
		memory[16'h5a09] <= 8'h3b;
		memory[16'h5a0a] <= 8'hd7;
		memory[16'h5a0b] <= 8'hc2;
		memory[16'h5a0c] <= 8'h35;
		memory[16'h5a0d] <= 8'h6a;
		memory[16'h5a0e] <= 8'h55;
		memory[16'h5a0f] <= 8'h1b;
		memory[16'h5a10] <= 8'h6a;
		memory[16'h5a11] <= 8'h41;
		memory[16'h5a12] <= 8'ha;
		memory[16'h5a13] <= 8'ha9;
		memory[16'h5a14] <= 8'hd2;
		memory[16'h5a15] <= 8'h42;
		memory[16'h5a16] <= 8'h66;
		memory[16'h5a17] <= 8'h86;
		memory[16'h5a18] <= 8'hd1;
		memory[16'h5a19] <= 8'hb6;
		memory[16'h5a1a] <= 8'h80;
		memory[16'h5a1b] <= 8'h3;
		memory[16'h5a1c] <= 8'h65;
		memory[16'h5a1d] <= 8'h94;
		memory[16'h5a1e] <= 8'h93;
		memory[16'h5a1f] <= 8'h19;
		memory[16'h5a20] <= 8'he5;
		memory[16'h5a21] <= 8'h39;
		memory[16'h5a22] <= 8'hd2;
		memory[16'h5a23] <= 8'haa;
		memory[16'h5a24] <= 8'h91;
		memory[16'h5a25] <= 8'hd8;
		memory[16'h5a26] <= 8'h11;
		memory[16'h5a27] <= 8'h6a;
		memory[16'h5a28] <= 8'h13;
		memory[16'h5a29] <= 8'he9;
		memory[16'h5a2a] <= 8'h2c;
		memory[16'h5a2b] <= 8'h48;
		memory[16'h5a2c] <= 8'h53;
		memory[16'h5a2d] <= 8'h81;
		memory[16'h5a2e] <= 8'h63;
		memory[16'h5a2f] <= 8'hbd;
		memory[16'h5a30] <= 8'hc3;
		memory[16'h5a31] <= 8'h6d;
		memory[16'h5a32] <= 8'h66;
		memory[16'h5a33] <= 8'h95;
		memory[16'h5a34] <= 8'haf;
		memory[16'h5a35] <= 8'hcd;
		memory[16'h5a36] <= 8'h1b;
		memory[16'h5a37] <= 8'h80;
		memory[16'h5a38] <= 8'h83;
		memory[16'h5a39] <= 8'h9b;
		memory[16'h5a3a] <= 8'h83;
		memory[16'h5a3b] <= 8'he8;
		memory[16'h5a3c] <= 8'h2f;
		memory[16'h5a3d] <= 8'h16;
		memory[16'h5a3e] <= 8'h1;
		memory[16'h5a3f] <= 8'h15;
		memory[16'h5a40] <= 8'h4f;
		memory[16'h5a41] <= 8'hd3;
		memory[16'h5a42] <= 8'hbf;
		memory[16'h5a43] <= 8'he1;
		memory[16'h5a44] <= 8'hab;
		memory[16'h5a45] <= 8'hd0;
		memory[16'h5a46] <= 8'h4b;
		memory[16'h5a47] <= 8'hbe;
		memory[16'h5a48] <= 8'hb9;
		memory[16'h5a49] <= 8'h77;
		memory[16'h5a4a] <= 8'h6;
		memory[16'h5a4b] <= 8'hc;
		memory[16'h5a4c] <= 8'hf8;
		memory[16'h5a4d] <= 8'h69;
		memory[16'h5a4e] <= 8'hc9;
		memory[16'h5a4f] <= 8'hbb;
		memory[16'h5a50] <= 8'hd6;
		memory[16'h5a51] <= 8'h30;
		memory[16'h5a52] <= 8'h50;
		memory[16'h5a53] <= 8'h85;
		memory[16'h5a54] <= 8'hfd;
		memory[16'h5a55] <= 8'h6b;
		memory[16'h5a56] <= 8'h5;
		memory[16'h5a57] <= 8'h80;
		memory[16'h5a58] <= 8'h6;
		memory[16'h5a59] <= 8'h89;
		memory[16'h5a5a] <= 8'h69;
		memory[16'h5a5b] <= 8'h36;
		memory[16'h5a5c] <= 8'h9f;
		memory[16'h5a5d] <= 8'h6a;
		memory[16'h5a5e] <= 8'h4b;
		memory[16'h5a5f] <= 8'hef;
		memory[16'h5a60] <= 8'h3e;
		memory[16'h5a61] <= 8'ha;
		memory[16'h5a62] <= 8'hd0;
		memory[16'h5a63] <= 8'he9;
		memory[16'h5a64] <= 8'hda;
		memory[16'h5a65] <= 8'h1b;
		memory[16'h5a66] <= 8'ha8;
		memory[16'h5a67] <= 8'h94;
		memory[16'h5a68] <= 8'h92;
		memory[16'h5a69] <= 8'hae;
		memory[16'h5a6a] <= 8'ha0;
		memory[16'h5a6b] <= 8'h8a;
		memory[16'h5a6c] <= 8'h18;
		memory[16'h5a6d] <= 8'h6a;
		memory[16'h5a6e] <= 8'h46;
		memory[16'h5a6f] <= 8'hee;
		memory[16'h5a70] <= 8'h9a;
		memory[16'h5a71] <= 8'h96;
		memory[16'h5a72] <= 8'h74;
		memory[16'h5a73] <= 8'h97;
		memory[16'h5a74] <= 8'h2;
		memory[16'h5a75] <= 8'h79;
		memory[16'h5a76] <= 8'h17;
		memory[16'h5a77] <= 8'h8;
		memory[16'h5a78] <= 8'h2;
		memory[16'h5a79] <= 8'h80;
		memory[16'h5a7a] <= 8'h3e;
		memory[16'h5a7b] <= 8'ha2;
		memory[16'h5a7c] <= 8'heb;
		memory[16'h5a7d] <= 8'h89;
		memory[16'h5a7e] <= 8'h91;
		memory[16'h5a7f] <= 8'h29;
		memory[16'h5a80] <= 8'h93;
		memory[16'h5a81] <= 8'h61;
		memory[16'h5a82] <= 8'h12;
		memory[16'h5a83] <= 8'h6e;
		memory[16'h5a84] <= 8'h7c;
		memory[16'h5a85] <= 8'hba;
		memory[16'h5a86] <= 8'h2;
		memory[16'h5a87] <= 8'he;
		memory[16'h5a88] <= 8'h69;
		memory[16'h5a89] <= 8'ha2;
		memory[16'h5a8a] <= 8'h98;
		memory[16'h5a8b] <= 8'h81;
		memory[16'h5a8c] <= 8'hc;
		memory[16'h5a8d] <= 8'hde;
		memory[16'h5a8e] <= 8'h6f;
		memory[16'h5a8f] <= 8'ha6;
		memory[16'h5a90] <= 8'h75;
		memory[16'h5a91] <= 8'he3;
		memory[16'h5a92] <= 8'h3d;
		memory[16'h5a93] <= 8'h77;
		memory[16'h5a94] <= 8'h5d;
		memory[16'h5a95] <= 8'h55;
		memory[16'h5a96] <= 8'h7f;
		memory[16'h5a97] <= 8'h5f;
		memory[16'h5a98] <= 8'hd5;
		memory[16'h5a99] <= 8'hbe;
		memory[16'h5a9a] <= 8'h1;
		memory[16'h5a9b] <= 8'hc0;
		memory[16'h5a9c] <= 8'h47;
		memory[16'h5a9d] <= 8'h92;
		memory[16'h5a9e] <= 8'he9;
		memory[16'h5a9f] <= 8'hdb;
		memory[16'h5aa0] <= 8'hf3;
		memory[16'h5aa1] <= 8'hfc;
		memory[16'h5aa2] <= 8'h49;
		memory[16'h5aa3] <= 8'h6f;
		memory[16'h5aa4] <= 8'hb6;
		memory[16'h5aa5] <= 8'h4b;
		memory[16'h5aa6] <= 8'h7d;
		memory[16'h5aa7] <= 8'h1f;
		memory[16'h5aa8] <= 8'hed;
		memory[16'h5aa9] <= 8'h16;
		memory[16'h5aaa] <= 8'ha0;
		memory[16'h5aab] <= 8'hfa;
		memory[16'h5aac] <= 8'hf4;
		memory[16'h5aad] <= 8'h10;
		memory[16'h5aae] <= 8'ha0;
		memory[16'h5aaf] <= 8'h69;
		memory[16'h5ab0] <= 8'hf3;
		memory[16'h5ab1] <= 8'hde;
		memory[16'h5ab2] <= 8'he0;
		memory[16'h5ab3] <= 8'h50;
		memory[16'h5ab4] <= 8'h33;
		memory[16'h5ab5] <= 8'h60;
		memory[16'h5ab6] <= 8'hb0;
		memory[16'h5ab7] <= 8'h8;
		memory[16'h5ab8] <= 8'h1e;
		memory[16'h5ab9] <= 8'hb1;
		memory[16'h5aba] <= 8'hc9;
		memory[16'h5abb] <= 8'h65;
		memory[16'h5abc] <= 8'h44;
		memory[16'h5abd] <= 8'hb2;
		memory[16'h5abe] <= 8'h40;
		memory[16'h5abf] <= 8'h37;
		memory[16'h5ac0] <= 8'hae;
		memory[16'h5ac1] <= 8'h89;
		memory[16'h5ac2] <= 8'ha7;
		memory[16'h5ac3] <= 8'h65;
		memory[16'h5ac4] <= 8'hd4;
		memory[16'h5ac5] <= 8'h24;
		memory[16'h5ac6] <= 8'h84;
		memory[16'h5ac7] <= 8'hc2;
		memory[16'h5ac8] <= 8'h3a;
		memory[16'h5ac9] <= 8'h25;
		memory[16'h5aca] <= 8'hbc;
		memory[16'h5acb] <= 8'h2f;
		memory[16'h5acc] <= 8'h35;
		memory[16'h5acd] <= 8'h5c;
		memory[16'h5ace] <= 8'h98;
		memory[16'h5acf] <= 8'h28;
		memory[16'h5ad0] <= 8'h3a;
		memory[16'h5ad1] <= 8'h79;
		memory[16'h5ad2] <= 8'h79;
		memory[16'h5ad3] <= 8'h6d;
		memory[16'h5ad4] <= 8'hd9;
		memory[16'h5ad5] <= 8'h29;
		memory[16'h5ad6] <= 8'h76;
		memory[16'h5ad7] <= 8'hf7;
		memory[16'h5ad8] <= 8'hda;
		memory[16'h5ad9] <= 8'h3f;
		memory[16'h5ada] <= 8'h5c;
		memory[16'h5adb] <= 8'h1e;
		memory[16'h5adc] <= 8'hf1;
		memory[16'h5add] <= 8'h9d;
		memory[16'h5ade] <= 8'h56;
		memory[16'h5adf] <= 8'ha0;
		memory[16'h5ae0] <= 8'h26;
		memory[16'h5ae1] <= 8'hfd;
		memory[16'h5ae2] <= 8'h5;
		memory[16'h5ae3] <= 8'hfb;
		memory[16'h5ae4] <= 8'h21;
		memory[16'h5ae5] <= 8'h89;
		memory[16'h5ae6] <= 8'hbd;
		memory[16'h5ae7] <= 8'h5c;
		memory[16'h5ae8] <= 8'hae;
		memory[16'h5ae9] <= 8'h79;
		memory[16'h5aea] <= 8'h8b;
		memory[16'h5aeb] <= 8'he3;
		memory[16'h5aec] <= 8'hd5;
		memory[16'h5aed] <= 8'h23;
		memory[16'h5aee] <= 8'hc;
		memory[16'h5aef] <= 8'h10;
		memory[16'h5af0] <= 8'h9c;
		memory[16'h5af1] <= 8'h85;
		memory[16'h5af2] <= 8'h7d;
		memory[16'h5af3] <= 8'h75;
		memory[16'h5af4] <= 8'hae;
		memory[16'h5af5] <= 8'hf3;
		memory[16'h5af6] <= 8'h6c;
		memory[16'h5af7] <= 8'h88;
		memory[16'h5af8] <= 8'h32;
		memory[16'h5af9] <= 8'hc9;
		memory[16'h5afa] <= 8'ha7;
		memory[16'h5afb] <= 8'h24;
		memory[16'h5afc] <= 8'h66;
		memory[16'h5afd] <= 8'hfd;
		memory[16'h5afe] <= 8'hc4;
		memory[16'h5aff] <= 8'h8c;
		memory[16'h5b00] <= 8'hfa;
		memory[16'h5b01] <= 8'hc9;
		memory[16'h5b02] <= 8'h87;
		memory[16'h5b03] <= 8'h1b;
		memory[16'h5b04] <= 8'h52;
		memory[16'h5b05] <= 8'h44;
		memory[16'h5b06] <= 8'h77;
		memory[16'h5b07] <= 8'h1;
		memory[16'h5b08] <= 8'hbd;
		memory[16'h5b09] <= 8'h2;
		memory[16'h5b0a] <= 8'he4;
		memory[16'h5b0b] <= 8'h93;
		memory[16'h5b0c] <= 8'h26;
		memory[16'h5b0d] <= 8'hf0;
		memory[16'h5b0e] <= 8'ha3;
		memory[16'h5b0f] <= 8'hc2;
		memory[16'h5b10] <= 8'h75;
		memory[16'h5b11] <= 8'h20;
		memory[16'h5b12] <= 8'h38;
		memory[16'h5b13] <= 8'h23;
		memory[16'h5b14] <= 8'h14;
		memory[16'h5b15] <= 8'ha4;
		memory[16'h5b16] <= 8'hac;
		memory[16'h5b17] <= 8'h46;
		memory[16'h5b18] <= 8'h6d;
		memory[16'h5b19] <= 8'h53;
		memory[16'h5b1a] <= 8'h6a;
		memory[16'h5b1b] <= 8'hd3;
		memory[16'h5b1c] <= 8'h50;
		memory[16'h5b1d] <= 8'h2e;
		memory[16'h5b1e] <= 8'h60;
		memory[16'h5b1f] <= 8'h4a;
		memory[16'h5b20] <= 8'hf7;
		memory[16'h5b21] <= 8'he7;
		memory[16'h5b22] <= 8'h65;
		memory[16'h5b23] <= 8'h4a;
		memory[16'h5b24] <= 8'h2c;
		memory[16'h5b25] <= 8'hdd;
		memory[16'h5b26] <= 8'h4b;
		memory[16'h5b27] <= 8'he9;
		memory[16'h5b28] <= 8'hdf;
		memory[16'h5b29] <= 8'h2f;
		memory[16'h5b2a] <= 8'h7c;
		memory[16'h5b2b] <= 8'h5;
		memory[16'h5b2c] <= 8'h20;
		memory[16'h5b2d] <= 8'h1f;
		memory[16'h5b2e] <= 8'hc8;
		memory[16'h5b2f] <= 8'h95;
		memory[16'h5b30] <= 8'h40;
		memory[16'h5b31] <= 8'h0;
		memory[16'h5b32] <= 8'hb9;
		memory[16'h5b33] <= 8'h54;
		memory[16'h5b34] <= 8'ha4;
		memory[16'h5b35] <= 8'h65;
		memory[16'h5b36] <= 8'h9a;
		memory[16'h5b37] <= 8'h12;
		memory[16'h5b38] <= 8'hb8;
		memory[16'h5b39] <= 8'h5;
		memory[16'h5b3a] <= 8'he5;
		memory[16'h5b3b] <= 8'h8;
		memory[16'h5b3c] <= 8'h33;
		memory[16'h5b3d] <= 8'h45;
		memory[16'h5b3e] <= 8'h52;
		memory[16'h5b3f] <= 8'h2b;
		memory[16'h5b40] <= 8'h2d;
		memory[16'h5b41] <= 8'hb7;
		memory[16'h5b42] <= 8'h75;
		memory[16'h5b43] <= 8'h59;
		memory[16'h5b44] <= 8'h94;
		memory[16'h5b45] <= 8'hc0;
		memory[16'h5b46] <= 8'h42;
		memory[16'h5b47] <= 8'h74;
		memory[16'h5b48] <= 8'hef;
		memory[16'h5b49] <= 8'hbf;
		memory[16'h5b4a] <= 8'h79;
		memory[16'h5b4b] <= 8'hf;
		memory[16'h5b4c] <= 8'hde;
		memory[16'h5b4d] <= 8'h41;
		memory[16'h5b4e] <= 8'ha5;
		memory[16'h5b4f] <= 8'h1e;
		memory[16'h5b50] <= 8'h41;
		memory[16'h5b51] <= 8'h5e;
		memory[16'h5b52] <= 8'h72;
		memory[16'h5b53] <= 8'he6;
		memory[16'h5b54] <= 8'hc3;
		memory[16'h5b55] <= 8'hd;
		memory[16'h5b56] <= 8'hf8;
		memory[16'h5b57] <= 8'h7b;
		memory[16'h5b58] <= 8'h12;
		memory[16'h5b59] <= 8'hdd;
		memory[16'h5b5a] <= 8'h83;
		memory[16'h5b5b] <= 8'h45;
		memory[16'h5b5c] <= 8'h23;
		memory[16'h5b5d] <= 8'hd5;
		memory[16'h5b5e] <= 8'h70;
		memory[16'h5b5f] <= 8'h50;
		memory[16'h5b60] <= 8'h8c;
		memory[16'h5b61] <= 8'he5;
		memory[16'h5b62] <= 8'ha9;
		memory[16'h5b63] <= 8'h21;
		memory[16'h5b64] <= 8'ha5;
		memory[16'h5b65] <= 8'heb;
		memory[16'h5b66] <= 8'h95;
		memory[16'h5b67] <= 8'h95;
		memory[16'h5b68] <= 8'haa;
		memory[16'h5b69] <= 8'he;
		memory[16'h5b6a] <= 8'ha4;
		memory[16'h5b6b] <= 8'h89;
		memory[16'h5b6c] <= 8'h50;
		memory[16'h5b6d] <= 8'h49;
		memory[16'h5b6e] <= 8'ha7;
		memory[16'h5b6f] <= 8'h91;
		memory[16'h5b70] <= 8'ha7;
		memory[16'h5b71] <= 8'h1a;
		memory[16'h5b72] <= 8'h77;
		memory[16'h5b73] <= 8'h6a;
		memory[16'h5b74] <= 8'h27;
		memory[16'h5b75] <= 8'h6f;
		memory[16'h5b76] <= 8'he5;
		memory[16'h5b77] <= 8'h39;
		memory[16'h5b78] <= 8'h4d;
		memory[16'h5b79] <= 8'h68;
		memory[16'h5b7a] <= 8'h7e;
		memory[16'h5b7b] <= 8'h70;
		memory[16'h5b7c] <= 8'h3d;
		memory[16'h5b7d] <= 8'hef;
		memory[16'h5b7e] <= 8'hc0;
		memory[16'h5b7f] <= 8'hca;
		memory[16'h5b80] <= 8'hd4;
		memory[16'h5b81] <= 8'h69;
		memory[16'h5b82] <= 8'heb;
		memory[16'h5b83] <= 8'h7a;
		memory[16'h5b84] <= 8'h54;
		memory[16'h5b85] <= 8'h80;
		memory[16'h5b86] <= 8'hf;
		memory[16'h5b87] <= 8'hff;
		memory[16'h5b88] <= 8'h8e;
		memory[16'h5b89] <= 8'hb3;
		memory[16'h5b8a] <= 8'h88;
		memory[16'h5b8b] <= 8'hde;
		memory[16'h5b8c] <= 8'hfd;
		memory[16'h5b8d] <= 8'h2f;
		memory[16'h5b8e] <= 8'h70;
		memory[16'h5b8f] <= 8'ha4;
		memory[16'h5b90] <= 8'h49;
		memory[16'h5b91] <= 8'he7;
		memory[16'h5b92] <= 8'hf;
		memory[16'h5b93] <= 8'h70;
		memory[16'h5b94] <= 8'h57;
		memory[16'h5b95] <= 8'hf4;
		memory[16'h5b96] <= 8'ha9;
		memory[16'h5b97] <= 8'ha4;
		memory[16'h5b98] <= 8'h5d;
		memory[16'h5b99] <= 8'h28;
		memory[16'h5b9a] <= 8'h14;
		memory[16'h5b9b] <= 8'h9a;
		memory[16'h5b9c] <= 8'h17;
		memory[16'h5b9d] <= 8'hd4;
		memory[16'h5b9e] <= 8'h64;
		memory[16'h5b9f] <= 8'heb;
		memory[16'h5ba0] <= 8'h3d;
		memory[16'h5ba1] <= 8'h4f;
		memory[16'h5ba2] <= 8'h65;
		memory[16'h5ba3] <= 8'h91;
		memory[16'h5ba4] <= 8'hcf;
		memory[16'h5ba5] <= 8'h74;
		memory[16'h5ba6] <= 8'h90;
		memory[16'h5ba7] <= 8'h5e;
		memory[16'h5ba8] <= 8'h28;
		memory[16'h5ba9] <= 8'h18;
		memory[16'h5baa] <= 8'h3c;
		memory[16'h5bab] <= 8'h25;
		memory[16'h5bac] <= 8'h48;
		memory[16'h5bad] <= 8'hac;
		memory[16'h5bae] <= 8'hc9;
		memory[16'h5baf] <= 8'h91;
		memory[16'h5bb0] <= 8'h94;
		memory[16'h5bb1] <= 8'hd8;
		memory[16'h5bb2] <= 8'h2;
		memory[16'h5bb3] <= 8'heb;
		memory[16'h5bb4] <= 8'hcd;
		memory[16'h5bb5] <= 8'hab;
		memory[16'h5bb6] <= 8'h8f;
		memory[16'h5bb7] <= 8'h2a;
		memory[16'h5bb8] <= 8'hd3;
		memory[16'h5bb9] <= 8'ha3;
		memory[16'h5bba] <= 8'hc4;
		memory[16'h5bbb] <= 8'hea;
		memory[16'h5bbc] <= 8'h77;
		memory[16'h5bbd] <= 8'h29;
		memory[16'h5bbe] <= 8'hd6;
		memory[16'h5bbf] <= 8'hb4;
		memory[16'h5bc0] <= 8'h78;
		memory[16'h5bc1] <= 8'h3b;
		memory[16'h5bc2] <= 8'h45;
		memory[16'h5bc3] <= 8'h48;
		memory[16'h5bc4] <= 8'hb0;
		memory[16'h5bc5] <= 8'hd6;
		memory[16'h5bc6] <= 8'ha6;
		memory[16'h5bc7] <= 8'hd8;
		memory[16'h5bc8] <= 8'hee;
		memory[16'h5bc9] <= 8'he2;
		memory[16'h5bca] <= 8'hfd;
		memory[16'h5bcb] <= 8'h36;
		memory[16'h5bcc] <= 8'h8f;
		memory[16'h5bcd] <= 8'hc6;
		memory[16'h5bce] <= 8'hc8;
		memory[16'h5bcf] <= 8'h23;
		memory[16'h5bd0] <= 8'h9f;
		memory[16'h5bd1] <= 8'hca;
		memory[16'h5bd2] <= 8'he;
		memory[16'h5bd3] <= 8'h6c;
		memory[16'h5bd4] <= 8'h75;
		memory[16'h5bd5] <= 8'h9d;
		memory[16'h5bd6] <= 8'h96;
		memory[16'h5bd7] <= 8'h49;
		memory[16'h5bd8] <= 8'h40;
		memory[16'h5bd9] <= 8'h5a;
		memory[16'h5bda] <= 8'h33;
		memory[16'h5bdb] <= 8'hb7;
		memory[16'h5bdc] <= 8'h83;
		memory[16'h5bdd] <= 8'h9;
		memory[16'h5bde] <= 8'h6b;
		memory[16'h5bdf] <= 8'hfc;
		memory[16'h5be0] <= 8'h45;
		memory[16'h5be1] <= 8'hb0;
		memory[16'h5be2] <= 8'h44;
		memory[16'h5be3] <= 8'hf5;
		memory[16'h5be4] <= 8'h86;
		memory[16'h5be5] <= 8'hea;
		memory[16'h5be6] <= 8'hcd;
		memory[16'h5be7] <= 8'h75;
		memory[16'h5be8] <= 8'hcc;
		memory[16'h5be9] <= 8'hca;
		memory[16'h5bea] <= 8'hab;
		memory[16'h5beb] <= 8'h5b;
		memory[16'h5bec] <= 8'h90;
		memory[16'h5bed] <= 8'h73;
		memory[16'h5bee] <= 8'h7e;
		memory[16'h5bef] <= 8'h2f;
		memory[16'h5bf0] <= 8'h3d;
		memory[16'h5bf1] <= 8'h8c;
		memory[16'h5bf2] <= 8'h9b;
		memory[16'h5bf3] <= 8'hb3;
		memory[16'h5bf4] <= 8'h29;
		memory[16'h5bf5] <= 8'h31;
		memory[16'h5bf6] <= 8'hfc;
		memory[16'h5bf7] <= 8'h69;
		memory[16'h5bf8] <= 8'h8c;
		memory[16'h5bf9] <= 8'h2f;
		memory[16'h5bfa] <= 8'h20;
		memory[16'h5bfb] <= 8'hf;
		memory[16'h5bfc] <= 8'h39;
		memory[16'h5bfd] <= 8'h8b;
		memory[16'h5bfe] <= 8'hb;
		memory[16'h5bff] <= 8'h7e;
		memory[16'h5c00] <= 8'h3c;
		memory[16'h5c01] <= 8'h4f;
		memory[16'h5c02] <= 8'h73;
		memory[16'h5c03] <= 8'hc2;
		memory[16'h5c04] <= 8'h39;
		memory[16'h5c05] <= 8'h40;
		memory[16'h5c06] <= 8'h37;
		memory[16'h5c07] <= 8'h6;
		memory[16'h5c08] <= 8'ha;
		memory[16'h5c09] <= 8'he3;
		memory[16'h5c0a] <= 8'h61;
		memory[16'h5c0b] <= 8'h9a;
		memory[16'h5c0c] <= 8'h56;
		memory[16'h5c0d] <= 8'he0;
		memory[16'h5c0e] <= 8'hca;
		memory[16'h5c0f] <= 8'h94;
		memory[16'h5c10] <= 8'h6c;
		memory[16'h5c11] <= 8'h65;
		memory[16'h5c12] <= 8'h47;
		memory[16'h5c13] <= 8'h96;
		memory[16'h5c14] <= 8'h97;
		memory[16'h5c15] <= 8'h43;
		memory[16'h5c16] <= 8'hff;
		memory[16'h5c17] <= 8'h23;
		memory[16'h5c18] <= 8'h72;
		memory[16'h5c19] <= 8'h20;
		memory[16'h5c1a] <= 8'h32;
		memory[16'h5c1b] <= 8'hab;
		memory[16'h5c1c] <= 8'hab;
		memory[16'h5c1d] <= 8'h3e;
		memory[16'h5c1e] <= 8'h29;
		memory[16'h5c1f] <= 8'he7;
		memory[16'h5c20] <= 8'h8d;
		memory[16'h5c21] <= 8'h9c;
		memory[16'h5c22] <= 8'haa;
		memory[16'h5c23] <= 8'hc7;
		memory[16'h5c24] <= 8'hdc;
		memory[16'h5c25] <= 8'he1;
		memory[16'h5c26] <= 8'hcd;
		memory[16'h5c27] <= 8'he6;
		memory[16'h5c28] <= 8'hc4;
		memory[16'h5c29] <= 8'h2e;
		memory[16'h5c2a] <= 8'h81;
		memory[16'h5c2b] <= 8'h1b;
		memory[16'h5c2c] <= 8'he;
		memory[16'h5c2d] <= 8'h4b;
		memory[16'h5c2e] <= 8'haf;
		memory[16'h5c2f] <= 8'h7b;
		memory[16'h5c30] <= 8'hb0;
		memory[16'h5c31] <= 8'hf6;
		memory[16'h5c32] <= 8'h11;
		memory[16'h5c33] <= 8'h47;
		memory[16'h5c34] <= 8'h39;
		memory[16'h5c35] <= 8'h10;
		memory[16'h5c36] <= 8'h6a;
		memory[16'h5c37] <= 8'hab;
		memory[16'h5c38] <= 8'h30;
		memory[16'h5c39] <= 8'h9d;
		memory[16'h5c3a] <= 8'h57;
		memory[16'h5c3b] <= 8'hdc;
		memory[16'h5c3c] <= 8'hdb;
		memory[16'h5c3d] <= 8'h80;
		memory[16'h5c3e] <= 8'hc3;
		memory[16'h5c3f] <= 8'h68;
		memory[16'h5c40] <= 8'h1d;
		memory[16'h5c41] <= 8'h6d;
		memory[16'h5c42] <= 8'h2f;
		memory[16'h5c43] <= 8'hf9;
		memory[16'h5c44] <= 8'h4f;
		memory[16'h5c45] <= 8'hfc;
		memory[16'h5c46] <= 8'he0;
		memory[16'h5c47] <= 8'h13;
		memory[16'h5c48] <= 8'h2b;
		memory[16'h5c49] <= 8'h61;
		memory[16'h5c4a] <= 8'h2e;
		memory[16'h5c4b] <= 8'h39;
		memory[16'h5c4c] <= 8'hac;
		memory[16'h5c4d] <= 8'hdd;
		memory[16'h5c4e] <= 8'hb4;
		memory[16'h5c4f] <= 8'h5c;
		memory[16'h5c50] <= 8'hd3;
		memory[16'h5c51] <= 8'hc5;
		memory[16'h5c52] <= 8'ha4;
		memory[16'h5c53] <= 8'hc;
		memory[16'h5c54] <= 8'hd6;
		memory[16'h5c55] <= 8'he;
		memory[16'h5c56] <= 8'hb8;
		memory[16'h5c57] <= 8'h6;
		memory[16'h5c58] <= 8'hab;
		memory[16'h5c59] <= 8'hf;
		memory[16'h5c5a] <= 8'he2;
		memory[16'h5c5b] <= 8'h86;
		memory[16'h5c5c] <= 8'h8f;
		memory[16'h5c5d] <= 8'ha6;
		memory[16'h5c5e] <= 8'hef;
		memory[16'h5c5f] <= 8'hac;
		memory[16'h5c60] <= 8'h13;
		memory[16'h5c61] <= 8'h1e;
		memory[16'h5c62] <= 8'ha6;
		memory[16'h5c63] <= 8'h62;
		memory[16'h5c64] <= 8'h1b;
		memory[16'h5c65] <= 8'h86;
		memory[16'h5c66] <= 8'h76;
		memory[16'h5c67] <= 8'h46;
		memory[16'h5c68] <= 8'he7;
		memory[16'h5c69] <= 8'ha4;
		memory[16'h5c6a] <= 8'h7f;
		memory[16'h5c6b] <= 8'h93;
		memory[16'h5c6c] <= 8'h82;
		memory[16'h5c6d] <= 8'h34;
		memory[16'h5c6e] <= 8'hef;
		memory[16'h5c6f] <= 8'h55;
		memory[16'h5c70] <= 8'hf9;
		memory[16'h5c71] <= 8'h93;
		memory[16'h5c72] <= 8'h62;
		memory[16'h5c73] <= 8'hcf;
		memory[16'h5c74] <= 8'ha2;
		memory[16'h5c75] <= 8'h1a;
		memory[16'h5c76] <= 8'hd6;
		memory[16'h5c77] <= 8'h4d;
		memory[16'h5c78] <= 8'h29;
		memory[16'h5c79] <= 8'hb8;
		memory[16'h5c7a] <= 8'hd4;
		memory[16'h5c7b] <= 8'hb8;
		memory[16'h5c7c] <= 8'h5e;
		memory[16'h5c7d] <= 8'hc3;
		memory[16'h5c7e] <= 8'h65;
		memory[16'h5c7f] <= 8'h72;
		memory[16'h5c80] <= 8'he1;
		memory[16'h5c81] <= 8'hb;
		memory[16'h5c82] <= 8'hd4;
		memory[16'h5c83] <= 8'hfc;
		memory[16'h5c84] <= 8'h91;
		memory[16'h5c85] <= 8'h4a;
		memory[16'h5c86] <= 8'h42;
		memory[16'h5c87] <= 8'h78;
		memory[16'h5c88] <= 8'hef;
		memory[16'h5c89] <= 8'hc2;
		memory[16'h5c8a] <= 8'hb;
		memory[16'h5c8b] <= 8'h71;
		memory[16'h5c8c] <= 8'hf6;
		memory[16'h5c8d] <= 8'hfa;
		memory[16'h5c8e] <= 8'hc6;
		memory[16'h5c8f] <= 8'hef;
		memory[16'h5c90] <= 8'h8e;
		memory[16'h5c91] <= 8'h28;
		memory[16'h5c92] <= 8'hbf;
		memory[16'h5c93] <= 8'h30;
		memory[16'h5c94] <= 8'h42;
		memory[16'h5c95] <= 8'h95;
		memory[16'h5c96] <= 8'h7d;
		memory[16'h5c97] <= 8'h6b;
		memory[16'h5c98] <= 8'h4d;
		memory[16'h5c99] <= 8'h51;
		memory[16'h5c9a] <= 8'h24;
		memory[16'h5c9b] <= 8'hac;
		memory[16'h5c9c] <= 8'h14;
		memory[16'h5c9d] <= 8'h89;
		memory[16'h5c9e] <= 8'h1e;
		memory[16'h5c9f] <= 8'hf6;
		memory[16'h5ca0] <= 8'h94;
		memory[16'h5ca1] <= 8'hf2;
		memory[16'h5ca2] <= 8'hf2;
		memory[16'h5ca3] <= 8'h25;
		memory[16'h5ca4] <= 8'h3d;
		memory[16'h5ca5] <= 8'h35;
		memory[16'h5ca6] <= 8'h9d;
		memory[16'h5ca7] <= 8'h2c;
		memory[16'h5ca8] <= 8'hf7;
		memory[16'h5ca9] <= 8'ha8;
		memory[16'h5caa] <= 8'h9d;
		memory[16'h5cab] <= 8'hed;
		memory[16'h5cac] <= 8'ha2;
		memory[16'h5cad] <= 8'h63;
		memory[16'h5cae] <= 8'hdc;
		memory[16'h5caf] <= 8'h30;
		memory[16'h5cb0] <= 8'h8c;
		memory[16'h5cb1] <= 8'h9b;
		memory[16'h5cb2] <= 8'h60;
		memory[16'h5cb3] <= 8'hce;
		memory[16'h5cb4] <= 8'h30;
		memory[16'h5cb5] <= 8'hde;
		memory[16'h5cb6] <= 8'h3a;
		memory[16'h5cb7] <= 8'h7e;
		memory[16'h5cb8] <= 8'h2f;
		memory[16'h5cb9] <= 8'h5e;
		memory[16'h5cba] <= 8'h2a;
		memory[16'h5cbb] <= 8'h44;
		memory[16'h5cbc] <= 8'he7;
		memory[16'h5cbd] <= 8'h48;
		memory[16'h5cbe] <= 8'h3a;
		memory[16'h5cbf] <= 8'h7b;
		memory[16'h5cc0] <= 8'h3a;
		memory[16'h5cc1] <= 8'h2c;
		memory[16'h5cc2] <= 8'ha0;
		memory[16'h5cc3] <= 8'h77;
		memory[16'h5cc4] <= 8'h61;
		memory[16'h5cc5] <= 8'h3d;
		memory[16'h5cc6] <= 8'ha3;
		memory[16'h5cc7] <= 8'h58;
		memory[16'h5cc8] <= 8'he5;
		memory[16'h5cc9] <= 8'h40;
		memory[16'h5cca] <= 8'h45;
		memory[16'h5ccb] <= 8'h87;
		memory[16'h5ccc] <= 8'ha4;
		memory[16'h5ccd] <= 8'h22;
		memory[16'h5cce] <= 8'hb8;
		memory[16'h5ccf] <= 8'h30;
		memory[16'h5cd0] <= 8'hbd;
		memory[16'h5cd1] <= 8'h18;
		memory[16'h5cd2] <= 8'hfe;
		memory[16'h5cd3] <= 8'hee;
		memory[16'h5cd4] <= 8'hf6;
		memory[16'h5cd5] <= 8'h38;
		memory[16'h5cd6] <= 8'h6c;
		memory[16'h5cd7] <= 8'h26;
		memory[16'h5cd8] <= 8'h96;
		memory[16'h5cd9] <= 8'h96;
		memory[16'h5cda] <= 8'h6a;
		memory[16'h5cdb] <= 8'h7d;
		memory[16'h5cdc] <= 8'hde;
		memory[16'h5cdd] <= 8'ha4;
		memory[16'h5cde] <= 8'hf8;
		memory[16'h5cdf] <= 8'h18;
		memory[16'h5ce0] <= 8'hd0;
		memory[16'h5ce1] <= 8'h98;
		memory[16'h5ce2] <= 8'h90;
		memory[16'h5ce3] <= 8'h32;
		memory[16'h5ce4] <= 8'hd5;
		memory[16'h5ce5] <= 8'h33;
		memory[16'h5ce6] <= 8'h8a;
		memory[16'h5ce7] <= 8'hba;
		memory[16'h5ce8] <= 8'h74;
		memory[16'h5ce9] <= 8'hd0;
		memory[16'h5cea] <= 8'h42;
		memory[16'h5ceb] <= 8'h18;
		memory[16'h5cec] <= 8'hf2;
		memory[16'h5ced] <= 8'hfa;
		memory[16'h5cee] <= 8'h48;
		memory[16'h5cef] <= 8'haf;
		memory[16'h5cf0] <= 8'h12;
		memory[16'h5cf1] <= 8'h46;
		memory[16'h5cf2] <= 8'h9d;
		memory[16'h5cf3] <= 8'h9;
		memory[16'h5cf4] <= 8'h7f;
		memory[16'h5cf5] <= 8'h9;
		memory[16'h5cf6] <= 8'h2f;
		memory[16'h5cf7] <= 8'h15;
		memory[16'h5cf8] <= 8'h9f;
		memory[16'h5cf9] <= 8'h99;
		memory[16'h5cfa] <= 8'h93;
		memory[16'h5cfb] <= 8'h7d;
		memory[16'h5cfc] <= 8'h3d;
		memory[16'h5cfd] <= 8'h8b;
		memory[16'h5cfe] <= 8'h96;
		memory[16'h5cff] <= 8'hd;
		memory[16'h5d00] <= 8'h24;
		memory[16'h5d01] <= 8'h26;
		memory[16'h5d02] <= 8'h3f;
		memory[16'h5d03] <= 8'hf9;
		memory[16'h5d04] <= 8'h59;
		memory[16'h5d05] <= 8'hca;
		memory[16'h5d06] <= 8'hb4;
		memory[16'h5d07] <= 8'hcd;
		memory[16'h5d08] <= 8'h9a;
		memory[16'h5d09] <= 8'hf6;
		memory[16'h5d0a] <= 8'he5;
		memory[16'h5d0b] <= 8'h8c;
		memory[16'h5d0c] <= 8'hf0;
		memory[16'h5d0d] <= 8'h2d;
		memory[16'h5d0e] <= 8'h3b;
		memory[16'h5d0f] <= 8'h2;
		memory[16'h5d10] <= 8'h74;
		memory[16'h5d11] <= 8'hd9;
		memory[16'h5d12] <= 8'hb;
		memory[16'h5d13] <= 8'hf3;
		memory[16'h5d14] <= 8'he2;
		memory[16'h5d15] <= 8'h3a;
		memory[16'h5d16] <= 8'h8;
		memory[16'h5d17] <= 8'h82;
		memory[16'h5d18] <= 8'hd3;
		memory[16'h5d19] <= 8'h9b;
		memory[16'h5d1a] <= 8'hff;
		memory[16'h5d1b] <= 8'h10;
		memory[16'h5d1c] <= 8'h27;
		memory[16'h5d1d] <= 8'h95;
		memory[16'h5d1e] <= 8'h1e;
		memory[16'h5d1f] <= 8'h4b;
		memory[16'h5d20] <= 8'hbb;
		memory[16'h5d21] <= 8'h5d;
		memory[16'h5d22] <= 8'h44;
		memory[16'h5d23] <= 8'h15;
		memory[16'h5d24] <= 8'h27;
		memory[16'h5d25] <= 8'hf8;
		memory[16'h5d26] <= 8'he2;
		memory[16'h5d27] <= 8'hc1;
		memory[16'h5d28] <= 8'hee;
		memory[16'h5d29] <= 8'hc8;
		memory[16'h5d2a] <= 8'h4d;
		memory[16'h5d2b] <= 8'hde;
		memory[16'h5d2c] <= 8'hf5;
		memory[16'h5d2d] <= 8'h89;
		memory[16'h5d2e] <= 8'he1;
		memory[16'h5d2f] <= 8'h69;
		memory[16'h5d30] <= 8'h62;
		memory[16'h5d31] <= 8'hec;
		memory[16'h5d32] <= 8'h5c;
		memory[16'h5d33] <= 8'h44;
		memory[16'h5d34] <= 8'h27;
		memory[16'h5d35] <= 8'h65;
		memory[16'h5d36] <= 8'hc6;
		memory[16'h5d37] <= 8'hfa;
		memory[16'h5d38] <= 8'h0;
		memory[16'h5d39] <= 8'hc6;
		memory[16'h5d3a] <= 8'hb;
		memory[16'h5d3b] <= 8'h27;
		memory[16'h5d3c] <= 8'h5b;
		memory[16'h5d3d] <= 8'h29;
		memory[16'h5d3e] <= 8'h72;
		memory[16'h5d3f] <= 8'h17;
		memory[16'h5d40] <= 8'h86;
		memory[16'h5d41] <= 8'hb7;
		memory[16'h5d42] <= 8'h2c;
		memory[16'h5d43] <= 8'hae;
		memory[16'h5d44] <= 8'haf;
		memory[16'h5d45] <= 8'he;
		memory[16'h5d46] <= 8'h6f;
		memory[16'h5d47] <= 8'h9e;
		memory[16'h5d48] <= 8'hd6;
		memory[16'h5d49] <= 8'hbd;
		memory[16'h5d4a] <= 8'h7c;
		memory[16'h5d4b] <= 8'hcc;
		memory[16'h5d4c] <= 8'h46;
		memory[16'h5d4d] <= 8'h5d;
		memory[16'h5d4e] <= 8'h35;
		memory[16'h5d4f] <= 8'ha8;
		memory[16'h5d50] <= 8'h4a;
		memory[16'h5d51] <= 8'h92;
		memory[16'h5d52] <= 8'hec;
		memory[16'h5d53] <= 8'h71;
		memory[16'h5d54] <= 8'hf7;
		memory[16'h5d55] <= 8'hb3;
		memory[16'h5d56] <= 8'h6b;
		memory[16'h5d57] <= 8'hf7;
		memory[16'h5d58] <= 8'h79;
		memory[16'h5d59] <= 8'h76;
		memory[16'h5d5a] <= 8'h1f;
		memory[16'h5d5b] <= 8'hd4;
		memory[16'h5d5c] <= 8'h9f;
		memory[16'h5d5d] <= 8'h91;
		memory[16'h5d5e] <= 8'heb;
		memory[16'h5d5f] <= 8'h26;
		memory[16'h5d60] <= 8'h48;
		memory[16'h5d61] <= 8'h17;
		memory[16'h5d62] <= 8'hd4;
		memory[16'h5d63] <= 8'hf8;
		memory[16'h5d64] <= 8'h26;
		memory[16'h5d65] <= 8'h43;
		memory[16'h5d66] <= 8'h96;
		memory[16'h5d67] <= 8'hfc;
		memory[16'h5d68] <= 8'h0;
		memory[16'h5d69] <= 8'h12;
		memory[16'h5d6a] <= 8'hc8;
		memory[16'h5d6b] <= 8'h46;
		memory[16'h5d6c] <= 8'h70;
		memory[16'h5d6d] <= 8'hfe;
		memory[16'h5d6e] <= 8'hee;
		memory[16'h5d6f] <= 8'hba;
		memory[16'h5d70] <= 8'h90;
		memory[16'h5d71] <= 8'hdb;
		memory[16'h5d72] <= 8'h2b;
		memory[16'h5d73] <= 8'h87;
		memory[16'h5d74] <= 8'h8e;
		memory[16'h5d75] <= 8'h96;
		memory[16'h5d76] <= 8'h7e;
		memory[16'h5d77] <= 8'h7;
		memory[16'h5d78] <= 8'hd;
		memory[16'h5d79] <= 8'h9d;
		memory[16'h5d7a] <= 8'hdb;
		memory[16'h5d7b] <= 8'hac;
		memory[16'h5d7c] <= 8'h2f;
		memory[16'h5d7d] <= 8'hc7;
		memory[16'h5d7e] <= 8'hd2;
		memory[16'h5d7f] <= 8'h77;
		memory[16'h5d80] <= 8'hde;
		memory[16'h5d81] <= 8'ha6;
		memory[16'h5d82] <= 8'h6f;
		memory[16'h5d83] <= 8'h4;
		memory[16'h5d84] <= 8'hea;
		memory[16'h5d85] <= 8'h5;
		memory[16'h5d86] <= 8'h1;
		memory[16'h5d87] <= 8'hea;
		memory[16'h5d88] <= 8'h18;
		memory[16'h5d89] <= 8'hc9;
		memory[16'h5d8a] <= 8'h31;
		memory[16'h5d8b] <= 8'h88;
		memory[16'h5d8c] <= 8'hc7;
		memory[16'h5d8d] <= 8'h1f;
		memory[16'h5d8e] <= 8'h42;
		memory[16'h5d8f] <= 8'h57;
		memory[16'h5d90] <= 8'hfa;
		memory[16'h5d91] <= 8'h6d;
		memory[16'h5d92] <= 8'hde;
		memory[16'h5d93] <= 8'h88;
		memory[16'h5d94] <= 8'h3;
		memory[16'h5d95] <= 8'h5d;
		memory[16'h5d96] <= 8'h8f;
		memory[16'h5d97] <= 8'h10;
		memory[16'h5d98] <= 8'hfa;
		memory[16'h5d99] <= 8'h6b;
		memory[16'h5d9a] <= 8'hbd;
		memory[16'h5d9b] <= 8'h29;
		memory[16'h5d9c] <= 8'h32;
		memory[16'h5d9d] <= 8'h8f;
		memory[16'h5d9e] <= 8'ha1;
		memory[16'h5d9f] <= 8'h10;
		memory[16'h5da0] <= 8'h36;
		memory[16'h5da1] <= 8'h10;
		memory[16'h5da2] <= 8'h15;
		memory[16'h5da3] <= 8'h20;
		memory[16'h5da4] <= 8'h16;
		memory[16'h5da5] <= 8'h16;
		memory[16'h5da6] <= 8'ha;
		memory[16'h5da7] <= 8'h2e;
		memory[16'h5da8] <= 8'hdf;
		memory[16'h5da9] <= 8'h3b;
		memory[16'h5daa] <= 8'hb6;
		memory[16'h5dab] <= 8'ha7;
		memory[16'h5dac] <= 8'h5b;
		memory[16'h5dad] <= 8'hf8;
		memory[16'h5dae] <= 8'hfe;
		memory[16'h5daf] <= 8'h55;
		memory[16'h5db0] <= 8'h65;
		memory[16'h5db1] <= 8'hdd;
		memory[16'h5db2] <= 8'hde;
		memory[16'h5db3] <= 8'h68;
		memory[16'h5db4] <= 8'h3a;
		memory[16'h5db5] <= 8'h6d;
		memory[16'h5db6] <= 8'h79;
		memory[16'h5db7] <= 8'h34;
		memory[16'h5db8] <= 8'hd8;
		memory[16'h5db9] <= 8'h36;
		memory[16'h5dba] <= 8'h5e;
		memory[16'h5dbb] <= 8'ha;
		memory[16'h5dbc] <= 8'hc5;
		memory[16'h5dbd] <= 8'hff;
		memory[16'h5dbe] <= 8'h1b;
		memory[16'h5dbf] <= 8'hfb;
		memory[16'h5dc0] <= 8'hf;
		memory[16'h5dc1] <= 8'h30;
		memory[16'h5dc2] <= 8'h1b;
		memory[16'h5dc3] <= 8'h25;
		memory[16'h5dc4] <= 8'h46;
		memory[16'h5dc5] <= 8'h26;
		memory[16'h5dc6] <= 8'h53;
		memory[16'h5dc7] <= 8'h25;
		memory[16'h5dc8] <= 8'h61;
		memory[16'h5dc9] <= 8'h9;
		memory[16'h5dca] <= 8'hcc;
		memory[16'h5dcb] <= 8'hbc;
		memory[16'h5dcc] <= 8'h1;
		memory[16'h5dcd] <= 8'hcb;
		memory[16'h5dce] <= 8'h12;
		memory[16'h5dcf] <= 8'h66;
		memory[16'h5dd0] <= 8'ha8;
		memory[16'h5dd1] <= 8'hf0;
		memory[16'h5dd2] <= 8'hcf;
		memory[16'h5dd3] <= 8'he2;
		memory[16'h5dd4] <= 8'h5d;
		memory[16'h5dd5] <= 8'h48;
		memory[16'h5dd6] <= 8'h16;
		memory[16'h5dd7] <= 8'h36;
		memory[16'h5dd8] <= 8'h7e;
		memory[16'h5dd9] <= 8'h74;
		memory[16'h5dda] <= 8'h40;
		memory[16'h5ddb] <= 8'h43;
		memory[16'h5ddc] <= 8'h73;
		memory[16'h5ddd] <= 8'h5b;
		memory[16'h5dde] <= 8'h3f;
		memory[16'h5ddf] <= 8'h83;
		memory[16'h5de0] <= 8'h8b;
		memory[16'h5de1] <= 8'h5a;
		memory[16'h5de2] <= 8'ha8;
		memory[16'h5de3] <= 8'hd1;
		memory[16'h5de4] <= 8'h80;
		memory[16'h5de5] <= 8'hfc;
		memory[16'h5de6] <= 8'hf7;
		memory[16'h5de7] <= 8'he2;
		memory[16'h5de8] <= 8'h5;
		memory[16'h5de9] <= 8'hc3;
		memory[16'h5dea] <= 8'h9e;
		memory[16'h5deb] <= 8'h7;
		memory[16'h5dec] <= 8'h8e;
		memory[16'h5ded] <= 8'hb0;
		memory[16'h5dee] <= 8'h6d;
		memory[16'h5def] <= 8'h36;
		memory[16'h5df0] <= 8'ha0;
		memory[16'h5df1] <= 8'h3c;
		memory[16'h5df2] <= 8'h18;
		memory[16'h5df3] <= 8'hfe;
		memory[16'h5df4] <= 8'h84;
		memory[16'h5df5] <= 8'h2f;
		memory[16'h5df6] <= 8'h34;
		memory[16'h5df7] <= 8'h2;
		memory[16'h5df8] <= 8'ha3;
		memory[16'h5df9] <= 8'h74;
		memory[16'h5dfa] <= 8'h46;
		memory[16'h5dfb] <= 8'h17;
		memory[16'h5dfc] <= 8'hd0;
		memory[16'h5dfd] <= 8'h85;
		memory[16'h5dfe] <= 8'h9a;
		memory[16'h5dff] <= 8'h5b;
		memory[16'h5e00] <= 8'hdf;
		memory[16'h5e01] <= 8'h42;
		memory[16'h5e02] <= 8'h2d;
		memory[16'h5e03] <= 8'h60;
		memory[16'h5e04] <= 8'h3e;
		memory[16'h5e05] <= 8'h24;
		memory[16'h5e06] <= 8'h42;
		memory[16'h5e07] <= 8'h44;
		memory[16'h5e08] <= 8'he7;
		memory[16'h5e09] <= 8'he0;
		memory[16'h5e0a] <= 8'h4b;
		memory[16'h5e0b] <= 8'h76;
		memory[16'h5e0c] <= 8'h91;
		memory[16'h5e0d] <= 8'hb8;
		memory[16'h5e0e] <= 8'hac;
		memory[16'h5e0f] <= 8'h31;
		memory[16'h5e10] <= 8'hf5;
		memory[16'h5e11] <= 8'hc5;
		memory[16'h5e12] <= 8'h2f;
		memory[16'h5e13] <= 8'h79;
		memory[16'h5e14] <= 8'hf4;
		memory[16'h5e15] <= 8'h63;
		memory[16'h5e16] <= 8'h7c;
		memory[16'h5e17] <= 8'h97;
		memory[16'h5e18] <= 8'hd8;
		memory[16'h5e19] <= 8'hc2;
		memory[16'h5e1a] <= 8'hae;
		memory[16'h5e1b] <= 8'ha8;
		memory[16'h5e1c] <= 8'h47;
		memory[16'h5e1d] <= 8'h48;
		memory[16'h5e1e] <= 8'h3;
		memory[16'h5e1f] <= 8'h26;
		memory[16'h5e20] <= 8'h8b;
		memory[16'h5e21] <= 8'h30;
		memory[16'h5e22] <= 8'h86;
		memory[16'h5e23] <= 8'hc9;
		memory[16'h5e24] <= 8'h54;
		memory[16'h5e25] <= 8'hc8;
		memory[16'h5e26] <= 8'hd;
		memory[16'h5e27] <= 8'h3c;
		memory[16'h5e28] <= 8'ha9;
		memory[16'h5e29] <= 8'h58;
		memory[16'h5e2a] <= 8'hb2;
		memory[16'h5e2b] <= 8'h3a;
		memory[16'h5e2c] <= 8'h11;
		memory[16'h5e2d] <= 8'h5e;
		memory[16'h5e2e] <= 8'h6b;
		memory[16'h5e2f] <= 8'h6;
		memory[16'h5e30] <= 8'h23;
		memory[16'h5e31] <= 8'h9b;
		memory[16'h5e32] <= 8'h7f;
		memory[16'h5e33] <= 8'h17;
		memory[16'h5e34] <= 8'hfe;
		memory[16'h5e35] <= 8'hfb;
		memory[16'h5e36] <= 8'haf;
		memory[16'h5e37] <= 8'hd6;
		memory[16'h5e38] <= 8'hbd;
		memory[16'h5e39] <= 8'h5d;
		memory[16'h5e3a] <= 8'h7e;
		memory[16'h5e3b] <= 8'h4;
		memory[16'h5e3c] <= 8'ha6;
		memory[16'h5e3d] <= 8'h82;
		memory[16'h5e3e] <= 8'h2b;
		memory[16'h5e3f] <= 8'h31;
		memory[16'h5e40] <= 8'hb2;
		memory[16'h5e41] <= 8'hb1;
		memory[16'h5e42] <= 8'hfa;
		memory[16'h5e43] <= 8'h7;
		memory[16'h5e44] <= 8'h7a;
		memory[16'h5e45] <= 8'h8;
		memory[16'h5e46] <= 8'h43;
		memory[16'h5e47] <= 8'h23;
		memory[16'h5e48] <= 8'h60;
		memory[16'h5e49] <= 8'hf5;
		memory[16'h5e4a] <= 8'h5d;
		memory[16'h5e4b] <= 8'h71;
		memory[16'h5e4c] <= 8'h53;
		memory[16'h5e4d] <= 8'hc8;
		memory[16'h5e4e] <= 8'h77;
		memory[16'h5e4f] <= 8'h77;
		memory[16'h5e50] <= 8'h63;
		memory[16'h5e51] <= 8'hf7;
		memory[16'h5e52] <= 8'h8e;
		memory[16'h5e53] <= 8'h62;
		memory[16'h5e54] <= 8'hf2;
		memory[16'h5e55] <= 8'h3d;
		memory[16'h5e56] <= 8'h38;
		memory[16'h5e57] <= 8'hb0;
		memory[16'h5e58] <= 8'h9b;
		memory[16'h5e59] <= 8'hb7;
		memory[16'h5e5a] <= 8'hb4;
		memory[16'h5e5b] <= 8'h41;
		memory[16'h5e5c] <= 8'h39;
		memory[16'h5e5d] <= 8'hdf;
		memory[16'h5e5e] <= 8'h72;
		memory[16'h5e5f] <= 8'heb;
		memory[16'h5e60] <= 8'h91;
		memory[16'h5e61] <= 8'h6c;
		memory[16'h5e62] <= 8'hf2;
		memory[16'h5e63] <= 8'hb;
		memory[16'h5e64] <= 8'h74;
		memory[16'h5e65] <= 8'h35;
		memory[16'h5e66] <= 8'h2e;
		memory[16'h5e67] <= 8'hd5;
		memory[16'h5e68] <= 8'h2a;
		memory[16'h5e69] <= 8'h8b;
		memory[16'h5e6a] <= 8'h46;
		memory[16'h5e6b] <= 8'h7e;
		memory[16'h5e6c] <= 8'h53;
		memory[16'h5e6d] <= 8'hbe;
		memory[16'h5e6e] <= 8'hf5;
		memory[16'h5e6f] <= 8'hb7;
		memory[16'h5e70] <= 8'hb5;
		memory[16'h5e71] <= 8'h83;
		memory[16'h5e72] <= 8'h19;
		memory[16'h5e73] <= 8'ha7;
		memory[16'h5e74] <= 8'hc1;
		memory[16'h5e75] <= 8'h51;
		memory[16'h5e76] <= 8'h57;
		memory[16'h5e77] <= 8'h5c;
		memory[16'h5e78] <= 8'h8;
		memory[16'h5e79] <= 8'hc;
		memory[16'h5e7a] <= 8'h9d;
		memory[16'h5e7b] <= 8'h41;
		memory[16'h5e7c] <= 8'heb;
		memory[16'h5e7d] <= 8'hf;
		memory[16'h5e7e] <= 8'h2d;
		memory[16'h5e7f] <= 8'h7c;
		memory[16'h5e80] <= 8'h7b;
		memory[16'h5e81] <= 8'h1f;
		memory[16'h5e82] <= 8'h87;
		memory[16'h5e83] <= 8'hf0;
		memory[16'h5e84] <= 8'h55;
		memory[16'h5e85] <= 8'hb5;
		memory[16'h5e86] <= 8'hc5;
		memory[16'h5e87] <= 8'h7f;
		memory[16'h5e88] <= 8'h40;
		memory[16'h5e89] <= 8'hb;
		memory[16'h5e8a] <= 8'hfd;
		memory[16'h5e8b] <= 8'h94;
		memory[16'h5e8c] <= 8'hc9;
		memory[16'h5e8d] <= 8'hf2;
		memory[16'h5e8e] <= 8'h4b;
		memory[16'h5e8f] <= 8'h7e;
		memory[16'h5e90] <= 8'h76;
		memory[16'h5e91] <= 8'h64;
		memory[16'h5e92] <= 8'h26;
		memory[16'h5e93] <= 8'h37;
		memory[16'h5e94] <= 8'hb5;
		memory[16'h5e95] <= 8'h7d;
		memory[16'h5e96] <= 8'h93;
		memory[16'h5e97] <= 8'hbe;
		memory[16'h5e98] <= 8'h89;
		memory[16'h5e99] <= 8'h30;
		memory[16'h5e9a] <= 8'hff;
		memory[16'h5e9b] <= 8'h75;
		memory[16'h5e9c] <= 8'h3f;
		memory[16'h5e9d] <= 8'h2c;
		memory[16'h5e9e] <= 8'hf1;
		memory[16'h5e9f] <= 8'hba;
		memory[16'h5ea0] <= 8'h4c;
		memory[16'h5ea1] <= 8'h79;
		memory[16'h5ea2] <= 8'haa;
		memory[16'h5ea3] <= 8'ha1;
		memory[16'h5ea4] <= 8'h2e;
		memory[16'h5ea5] <= 8'h6f;
		memory[16'h5ea6] <= 8'h20;
		memory[16'h5ea7] <= 8'h6f;
		memory[16'h5ea8] <= 8'h7b;
		memory[16'h5ea9] <= 8'h1e;
		memory[16'h5eaa] <= 8'h3;
		memory[16'h5eab] <= 8'h44;
		memory[16'h5eac] <= 8'h10;
		memory[16'h5ead] <= 8'h4e;
		memory[16'h5eae] <= 8'hc3;
		memory[16'h5eaf] <= 8'h86;
		memory[16'h5eb0] <= 8'hb2;
		memory[16'h5eb1] <= 8'he9;
		memory[16'h5eb2] <= 8'hbd;
		memory[16'h5eb3] <= 8'h67;
		memory[16'h5eb4] <= 8'h66;
		memory[16'h5eb5] <= 8'h50;
		memory[16'h5eb6] <= 8'h25;
		memory[16'h5eb7] <= 8'hf0;
		memory[16'h5eb8] <= 8'h80;
		memory[16'h5eb9] <= 8'h25;
		memory[16'h5eba] <= 8'h65;
		memory[16'h5ebb] <= 8'hbf;
		memory[16'h5ebc] <= 8'h51;
		memory[16'h5ebd] <= 8'h56;
		memory[16'h5ebe] <= 8'h7a;
		memory[16'h5ebf] <= 8'h9d;
		memory[16'h5ec0] <= 8'hcf;
		memory[16'h5ec1] <= 8'h24;
		memory[16'h5ec2] <= 8'h3e;
		memory[16'h5ec3] <= 8'hfe;
		memory[16'h5ec4] <= 8'h94;
		memory[16'h5ec5] <= 8'h5f;
		memory[16'h5ec6] <= 8'h6d;
		memory[16'h5ec7] <= 8'hf;
		memory[16'h5ec8] <= 8'h7d;
		memory[16'h5ec9] <= 8'h70;
		memory[16'h5eca] <= 8'h53;
		memory[16'h5ecb] <= 8'h8d;
		memory[16'h5ecc] <= 8'hbe;
		memory[16'h5ecd] <= 8'h16;
		memory[16'h5ece] <= 8'h14;
		memory[16'h5ecf] <= 8'h70;
		memory[16'h5ed0] <= 8'hff;
		memory[16'h5ed1] <= 8'hd1;
		memory[16'h5ed2] <= 8'hd7;
		memory[16'h5ed3] <= 8'h66;
		memory[16'h5ed4] <= 8'h22;
		memory[16'h5ed5] <= 8'hfd;
		memory[16'h5ed6] <= 8'h56;
		memory[16'h5ed7] <= 8'ha2;
		memory[16'h5ed8] <= 8'h22;
		memory[16'h5ed9] <= 8'hbb;
		memory[16'h5eda] <= 8'h62;
		memory[16'h5edb] <= 8'h73;
		memory[16'h5edc] <= 8'h11;
		memory[16'h5edd] <= 8'hdc;
		memory[16'h5ede] <= 8'h11;
		memory[16'h5edf] <= 8'he1;
		memory[16'h5ee0] <= 8'h0;
		memory[16'h5ee1] <= 8'h4f;
		memory[16'h5ee2] <= 8'hdf;
		memory[16'h5ee3] <= 8'h94;
		memory[16'h5ee4] <= 8'hae;
		memory[16'h5ee5] <= 8'h4c;
		memory[16'h5ee6] <= 8'ha3;
		memory[16'h5ee7] <= 8'h2b;
		memory[16'h5ee8] <= 8'hbc;
		memory[16'h5ee9] <= 8'hf7;
		memory[16'h5eea] <= 8'hb9;
		memory[16'h5eeb] <= 8'h7a;
		memory[16'h5eec] <= 8'hd;
		memory[16'h5eed] <= 8'hcd;
		memory[16'h5eee] <= 8'hea;
		memory[16'h5eef] <= 8'hd;
		memory[16'h5ef0] <= 8'h9e;
		memory[16'h5ef1] <= 8'hc1;
		memory[16'h5ef2] <= 8'h73;
		memory[16'h5ef3] <= 8'hc0;
		memory[16'h5ef4] <= 8'hbe;
		memory[16'h5ef5] <= 8'hc9;
		memory[16'h5ef6] <= 8'h63;
		memory[16'h5ef7] <= 8'he0;
		memory[16'h5ef8] <= 8'h84;
		memory[16'h5ef9] <= 8'hc5;
		memory[16'h5efa] <= 8'h54;
		memory[16'h5efb] <= 8'h95;
		memory[16'h5efc] <= 8'ha1;
		memory[16'h5efd] <= 8'h65;
		memory[16'h5efe] <= 8'h76;
		memory[16'h5eff] <= 8'ha1;
		memory[16'h5f00] <= 8'hb4;
		memory[16'h5f01] <= 8'h55;
		memory[16'h5f02] <= 8'h36;
		memory[16'h5f03] <= 8'h63;
		memory[16'h5f04] <= 8'ha1;
		memory[16'h5f05] <= 8'hd9;
		memory[16'h5f06] <= 8'h8e;
		memory[16'h5f07] <= 8'h5d;
		memory[16'h5f08] <= 8'hd0;
		memory[16'h5f09] <= 8'h47;
		memory[16'h5f0a] <= 8'hd7;
		memory[16'h5f0b] <= 8'hde;
		memory[16'h5f0c] <= 8'h14;
		memory[16'h5f0d] <= 8'hc1;
		memory[16'h5f0e] <= 8'heb;
		memory[16'h5f0f] <= 8'hb3;
		memory[16'h5f10] <= 8'h83;
		memory[16'h5f11] <= 8'h5e;
		memory[16'h5f12] <= 8'h73;
		memory[16'h5f13] <= 8'h41;
		memory[16'h5f14] <= 8'h27;
		memory[16'h5f15] <= 8'hd6;
		memory[16'h5f16] <= 8'h22;
		memory[16'h5f17] <= 8'hab;
		memory[16'h5f18] <= 8'h9b;
		memory[16'h5f19] <= 8'h76;
		memory[16'h5f1a] <= 8'h40;
		memory[16'h5f1b] <= 8'h3c;
		memory[16'h5f1c] <= 8'hdb;
		memory[16'h5f1d] <= 8'hb7;
		memory[16'h5f1e] <= 8'hde;
		memory[16'h5f1f] <= 8'h8f;
		memory[16'h5f20] <= 8'hc;
		memory[16'h5f21] <= 8'h14;
		memory[16'h5f22] <= 8'hf2;
		memory[16'h5f23] <= 8'hae;
		memory[16'h5f24] <= 8'hed;
		memory[16'h5f25] <= 8'h81;
		memory[16'h5f26] <= 8'hb;
		memory[16'h5f27] <= 8'hbe;
		memory[16'h5f28] <= 8'hc8;
		memory[16'h5f29] <= 8'he3;
		memory[16'h5f2a] <= 8'h9c;
		memory[16'h5f2b] <= 8'hdd;
		memory[16'h5f2c] <= 8'ha4;
		memory[16'h5f2d] <= 8'h87;
		memory[16'h5f2e] <= 8'h90;
		memory[16'h5f2f] <= 8'h27;
		memory[16'h5f30] <= 8'he5;
		memory[16'h5f31] <= 8'h3;
		memory[16'h5f32] <= 8'h69;
		memory[16'h5f33] <= 8'hc;
		memory[16'h5f34] <= 8'hda;
		memory[16'h5f35] <= 8'h8b;
		memory[16'h5f36] <= 8'hb7;
		memory[16'h5f37] <= 8'h75;
		memory[16'h5f38] <= 8'h1;
		memory[16'h5f39] <= 8'hf7;
		memory[16'h5f3a] <= 8'hb2;
		memory[16'h5f3b] <= 8'hdc;
		memory[16'h5f3c] <= 8'hae;
		memory[16'h5f3d] <= 8'h90;
		memory[16'h5f3e] <= 8'h6b;
		memory[16'h5f3f] <= 8'hbb;
		memory[16'h5f40] <= 8'ha4;
		memory[16'h5f41] <= 8'h5e;
		memory[16'h5f42] <= 8'h69;
		memory[16'h5f43] <= 8'h91;
		memory[16'h5f44] <= 8'hdf;
		memory[16'h5f45] <= 8'h74;
		memory[16'h5f46] <= 8'h4f;
		memory[16'h5f47] <= 8'ha7;
		memory[16'h5f48] <= 8'h57;
		memory[16'h5f49] <= 8'heb;
		memory[16'h5f4a] <= 8'h84;
		memory[16'h5f4b] <= 8'hfc;
		memory[16'h5f4c] <= 8'h72;
		memory[16'h5f4d] <= 8'h14;
		memory[16'h5f4e] <= 8'h23;
		memory[16'h5f4f] <= 8'h57;
		memory[16'h5f50] <= 8'h18;
		memory[16'h5f51] <= 8'h8c;
		memory[16'h5f52] <= 8'h63;
		memory[16'h5f53] <= 8'hf2;
		memory[16'h5f54] <= 8'h17;
		memory[16'h5f55] <= 8'h1a;
		memory[16'h5f56] <= 8'h67;
		memory[16'h5f57] <= 8'h18;
		memory[16'h5f58] <= 8'h12;
		memory[16'h5f59] <= 8'h19;
		memory[16'h5f5a] <= 8'hf4;
		memory[16'h5f5b] <= 8'hc0;
		memory[16'h5f5c] <= 8'ha9;
		memory[16'h5f5d] <= 8'h60;
		memory[16'h5f5e] <= 8'h7b;
		memory[16'h5f5f] <= 8'h4d;
		memory[16'h5f60] <= 8'hbe;
		memory[16'h5f61] <= 8'he4;
		memory[16'h5f62] <= 8'hdf;
		memory[16'h5f63] <= 8'h9d;
		memory[16'h5f64] <= 8'h59;
		memory[16'h5f65] <= 8'h2e;
		memory[16'h5f66] <= 8'h44;
		memory[16'h5f67] <= 8'hb0;
		memory[16'h5f68] <= 8'h1a;
		memory[16'h5f69] <= 8'hc9;
		memory[16'h5f6a] <= 8'hac;
		memory[16'h5f6b] <= 8'h8c;
		memory[16'h5f6c] <= 8'hdd;
		memory[16'h5f6d] <= 8'hd0;
		memory[16'h5f6e] <= 8'he4;
		memory[16'h5f6f] <= 8'hf5;
		memory[16'h5f70] <= 8'h5c;
		memory[16'h5f71] <= 8'h47;
		memory[16'h5f72] <= 8'he7;
		memory[16'h5f73] <= 8'h74;
		memory[16'h5f74] <= 8'h62;
		memory[16'h5f75] <= 8'h4f;
		memory[16'h5f76] <= 8'h8c;
		memory[16'h5f77] <= 8'h74;
		memory[16'h5f78] <= 8'h68;
		memory[16'h5f79] <= 8'h81;
		memory[16'h5f7a] <= 8'h34;
		memory[16'h5f7b] <= 8'h12;
		memory[16'h5f7c] <= 8'he1;
		memory[16'h5f7d] <= 8'hb0;
		memory[16'h5f7e] <= 8'h5f;
		memory[16'h5f7f] <= 8'h9f;
		memory[16'h5f80] <= 8'h94;
		memory[16'h5f81] <= 8'h3e;
		memory[16'h5f82] <= 8'h3c;
		memory[16'h5f83] <= 8'hed;
		memory[16'h5f84] <= 8'h6d;
		memory[16'h5f85] <= 8'h80;
		memory[16'h5f86] <= 8'h9e;
		memory[16'h5f87] <= 8'h87;
		memory[16'h5f88] <= 8'h49;
		memory[16'h5f89] <= 8'h4a;
		memory[16'h5f8a] <= 8'h13;
		memory[16'h5f8b] <= 8'h27;
		memory[16'h5f8c] <= 8'h1a;
		memory[16'h5f8d] <= 8'hf7;
		memory[16'h5f8e] <= 8'h1c;
		memory[16'h5f8f] <= 8'h77;
		memory[16'h5f90] <= 8'h3f;
		memory[16'h5f91] <= 8'h4;
		memory[16'h5f92] <= 8'heb;
		memory[16'h5f93] <= 8'ha1;
		memory[16'h5f94] <= 8'h53;
		memory[16'h5f95] <= 8'h77;
		memory[16'h5f96] <= 8'h15;
		memory[16'h5f97] <= 8'hbb;
		memory[16'h5f98] <= 8'hf8;
		memory[16'h5f99] <= 8'h49;
		memory[16'h5f9a] <= 8'hcd;
		memory[16'h5f9b] <= 8'hd9;
		memory[16'h5f9c] <= 8'hf9;
		memory[16'h5f9d] <= 8'h2d;
		memory[16'h5f9e] <= 8'h78;
		memory[16'h5f9f] <= 8'h8e;
		memory[16'h5fa0] <= 8'h6b;
		memory[16'h5fa1] <= 8'hb4;
		memory[16'h5fa2] <= 8'h7b;
		memory[16'h5fa3] <= 8'hd8;
		memory[16'h5fa4] <= 8'h35;
		memory[16'h5fa5] <= 8'h19;
		memory[16'h5fa6] <= 8'h5f;
		memory[16'h5fa7] <= 8'h7e;
		memory[16'h5fa8] <= 8'h64;
		memory[16'h5fa9] <= 8'h73;
		memory[16'h5faa] <= 8'ha5;
		memory[16'h5fab] <= 8'h7e;
		memory[16'h5fac] <= 8'h6a;
		memory[16'h5fad] <= 8'hc2;
		memory[16'h5fae] <= 8'hf5;
		memory[16'h5faf] <= 8'ha9;
		memory[16'h5fb0] <= 8'hc6;
		memory[16'h5fb1] <= 8'he0;
		memory[16'h5fb2] <= 8'h4a;
		memory[16'h5fb3] <= 8'h19;
		memory[16'h5fb4] <= 8'h58;
		memory[16'h5fb5] <= 8'h5f;
		memory[16'h5fb6] <= 8'hd4;
		memory[16'h5fb7] <= 8'h50;
		memory[16'h5fb8] <= 8'ha9;
		memory[16'h5fb9] <= 8'ha2;
		memory[16'h5fba] <= 8'h2a;
		memory[16'h5fbb] <= 8'ha2;
		memory[16'h5fbc] <= 8'hcf;
		memory[16'h5fbd] <= 8'ha2;
		memory[16'h5fbe] <= 8'h30;
		memory[16'h5fbf] <= 8'h3a;
		memory[16'h5fc0] <= 8'h57;
		memory[16'h5fc1] <= 8'hac;
		memory[16'h5fc2] <= 8'h13;
		memory[16'h5fc3] <= 8'h8c;
		memory[16'h5fc4] <= 8'hc5;
		memory[16'h5fc5] <= 8'h72;
		memory[16'h5fc6] <= 8'ha;
		memory[16'h5fc7] <= 8'h29;
		memory[16'h5fc8] <= 8'he5;
		memory[16'h5fc9] <= 8'hb0;
		memory[16'h5fca] <= 8'ha8;
		memory[16'h5fcb] <= 8'h50;
		memory[16'h5fcc] <= 8'h72;
		memory[16'h5fcd] <= 8'h9d;
		memory[16'h5fce] <= 8'hf9;
		memory[16'h5fcf] <= 8'h38;
		memory[16'h5fd0] <= 8'h7e;
		memory[16'h5fd1] <= 8'h44;
		memory[16'h5fd2] <= 8'h51;
		memory[16'h5fd3] <= 8'hd6;
		memory[16'h5fd4] <= 8'ha3;
		memory[16'h5fd5] <= 8'h25;
		memory[16'h5fd6] <= 8'h26;
		memory[16'h5fd7] <= 8'h4c;
		memory[16'h5fd8] <= 8'hc7;
		memory[16'h5fd9] <= 8'h50;
		memory[16'h5fda] <= 8'hef;
		memory[16'h5fdb] <= 8'h96;
		memory[16'h5fdc] <= 8'hf3;
		memory[16'h5fdd] <= 8'h1f;
		memory[16'h5fde] <= 8'hd1;
		memory[16'h5fdf] <= 8'h4a;
		memory[16'h5fe0] <= 8'hcb;
		memory[16'h5fe1] <= 8'he4;
		memory[16'h5fe2] <= 8'hd6;
		memory[16'h5fe3] <= 8'h91;
		memory[16'h5fe4] <= 8'h56;
		memory[16'h5fe5] <= 8'he0;
		memory[16'h5fe6] <= 8'hba;
		memory[16'h5fe7] <= 8'h3c;
		memory[16'h5fe8] <= 8'h90;
		memory[16'h5fe9] <= 8'h62;
		memory[16'h5fea] <= 8'h8c;
		memory[16'h5feb] <= 8'h2;
		memory[16'h5fec] <= 8'h0;
		memory[16'h5fed] <= 8'h85;
		memory[16'h5fee] <= 8'h3a;
		memory[16'h5fef] <= 8'h7e;
		memory[16'h5ff0] <= 8'hc9;
		memory[16'h5ff1] <= 8'h8b;
		memory[16'h5ff2] <= 8'h54;
		memory[16'h5ff3] <= 8'h6d;
		memory[16'h5ff4] <= 8'hb1;
		memory[16'h5ff5] <= 8'h7a;
		memory[16'h5ff6] <= 8'hb9;
		memory[16'h5ff7] <= 8'h78;
		memory[16'h5ff8] <= 8'hcb;
		memory[16'h5ff9] <= 8'ha8;
		memory[16'h5ffa] <= 8'hf;
		memory[16'h5ffb] <= 8'hbe;
		memory[16'h5ffc] <= 8'hc8;
		memory[16'h5ffd] <= 8'he0;
		memory[16'h5ffe] <= 8'h8;
		memory[16'h5fff] <= 8'h93;
		memory[16'h6000] <= 8'hc4;
		memory[16'h6001] <= 8'hde;
		memory[16'h6002] <= 8'h24;
		memory[16'h6003] <= 8'h1a;
		memory[16'h6004] <= 8'hbe;
		memory[16'h6005] <= 8'hdf;
		memory[16'h6006] <= 8'h56;
		memory[16'h6007] <= 8'h4f;
		memory[16'h6008] <= 8'h41;
		memory[16'h6009] <= 8'he2;
		memory[16'h600a] <= 8'h51;
		memory[16'h600b] <= 8'h41;
		memory[16'h600c] <= 8'h68;
		memory[16'h600d] <= 8'h8c;
		memory[16'h600e] <= 8'hbf;
		memory[16'h600f] <= 8'h31;
		memory[16'h6010] <= 8'h17;
		memory[16'h6011] <= 8'h13;
		memory[16'h6012] <= 8'h9e;
		memory[16'h6013] <= 8'hc8;
		memory[16'h6014] <= 8'h8e;
		memory[16'h6015] <= 8'h58;
		memory[16'h6016] <= 8'h41;
		memory[16'h6017] <= 8'h59;
		memory[16'h6018] <= 8'h0;
		memory[16'h6019] <= 8'h50;
		memory[16'h601a] <= 8'h17;
		memory[16'h601b] <= 8'hc8;
		memory[16'h601c] <= 8'h30;
		memory[16'h601d] <= 8'h1f;
		memory[16'h601e] <= 8'h5c;
		memory[16'h601f] <= 8'hf4;
		memory[16'h6020] <= 8'hfd;
		memory[16'h6021] <= 8'h80;
		memory[16'h6022] <= 8'he;
		memory[16'h6023] <= 8'hbb;
		memory[16'h6024] <= 8'h5f;
		memory[16'h6025] <= 8'h65;
		memory[16'h6026] <= 8'ha;
		memory[16'h6027] <= 8'ha1;
		memory[16'h6028] <= 8'h47;
		memory[16'h6029] <= 8'h5c;
		memory[16'h602a] <= 8'he2;
		memory[16'h602b] <= 8'haf;
		memory[16'h602c] <= 8'he8;
		memory[16'h602d] <= 8'ha2;
		memory[16'h602e] <= 8'he1;
		memory[16'h602f] <= 8'hff;
		memory[16'h6030] <= 8'hb5;
		memory[16'h6031] <= 8'h7f;
		memory[16'h6032] <= 8'hc8;
		memory[16'h6033] <= 8'h43;
		memory[16'h6034] <= 8'hd7;
		memory[16'h6035] <= 8'h9;
		memory[16'h6036] <= 8'h9c;
		memory[16'h6037] <= 8'hd8;
		memory[16'h6038] <= 8'h59;
		memory[16'h6039] <= 8'hb3;
		memory[16'h603a] <= 8'ha0;
		memory[16'h603b] <= 8'h89;
		memory[16'h603c] <= 8'hd2;
		memory[16'h603d] <= 8'hfc;
		memory[16'h603e] <= 8'h7d;
		memory[16'h603f] <= 8'hcf;
		memory[16'h6040] <= 8'h7d;
		memory[16'h6041] <= 8'h8b;
		memory[16'h6042] <= 8'h8b;
		memory[16'h6043] <= 8'hdc;
		memory[16'h6044] <= 8'hf0;
		memory[16'h6045] <= 8'h95;
		memory[16'h6046] <= 8'h7d;
		memory[16'h6047] <= 8'h38;
		memory[16'h6048] <= 8'hf1;
		memory[16'h6049] <= 8'h60;
		memory[16'h604a] <= 8'he7;
		memory[16'h604b] <= 8'hd9;
		memory[16'h604c] <= 8'h2;
		memory[16'h604d] <= 8'hc8;
		memory[16'h604e] <= 8'hd9;
		memory[16'h604f] <= 8'hb7;
		memory[16'h6050] <= 8'h48;
		memory[16'h6051] <= 8'ha1;
		memory[16'h6052] <= 8'hfb;
		memory[16'h6053] <= 8'h1f;
		memory[16'h6054] <= 8'haa;
		memory[16'h6055] <= 8'h97;
		memory[16'h6056] <= 8'hf7;
		memory[16'h6057] <= 8'h3;
		memory[16'h6058] <= 8'h4b;
		memory[16'h6059] <= 8'h98;
		memory[16'h605a] <= 8'h8c;
		memory[16'h605b] <= 8'h1d;
		memory[16'h605c] <= 8'h94;
		memory[16'h605d] <= 8'h9;
		memory[16'h605e] <= 8'hed;
		memory[16'h605f] <= 8'h11;
		memory[16'h6060] <= 8'h94;
		memory[16'h6061] <= 8'h78;
		memory[16'h6062] <= 8'hee;
		memory[16'h6063] <= 8'h85;
		memory[16'h6064] <= 8'hd;
		memory[16'h6065] <= 8'h6b;
		memory[16'h6066] <= 8'hbd;
		memory[16'h6067] <= 8'hff;
		memory[16'h6068] <= 8'hcb;
		memory[16'h6069] <= 8'ha4;
		memory[16'h606a] <= 8'hd8;
		memory[16'h606b] <= 8'hcd;
		memory[16'h606c] <= 8'h6d;
		memory[16'h606d] <= 8'hb1;
		memory[16'h606e] <= 8'h85;
		memory[16'h606f] <= 8'hb5;
		memory[16'h6070] <= 8'h52;
		memory[16'h6071] <= 8'h80;
		memory[16'h6072] <= 8'hd4;
		memory[16'h6073] <= 8'hfc;
		memory[16'h6074] <= 8'h17;
		memory[16'h6075] <= 8'hcc;
		memory[16'h6076] <= 8'hff;
		memory[16'h6077] <= 8'h62;
		memory[16'h6078] <= 8'h64;
		memory[16'h6079] <= 8'h8b;
		memory[16'h607a] <= 8'h80;
		memory[16'h607b] <= 8'hf8;
		memory[16'h607c] <= 8'h94;
		memory[16'h607d] <= 8'h6d;
		memory[16'h607e] <= 8'ha;
		memory[16'h607f] <= 8'h29;
		memory[16'h6080] <= 8'he5;
		memory[16'h6081] <= 8'hf8;
		memory[16'h6082] <= 8'hae;
		memory[16'h6083] <= 8'hf2;
		memory[16'h6084] <= 8'h63;
		memory[16'h6085] <= 8'h6b;
		memory[16'h6086] <= 8'hf1;
		memory[16'h6087] <= 8'h2f;
		memory[16'h6088] <= 8'hf;
		memory[16'h6089] <= 8'hca;
		memory[16'h608a] <= 8'hfc;
		memory[16'h608b] <= 8'h7c;
		memory[16'h608c] <= 8'h7b;
		memory[16'h608d] <= 8'h81;
		memory[16'h608e] <= 8'h31;
		memory[16'h608f] <= 8'hce;
		memory[16'h6090] <= 8'h1;
		memory[16'h6091] <= 8'h6;
		memory[16'h6092] <= 8'hca;
		memory[16'h6093] <= 8'h19;
		memory[16'h6094] <= 8'hd2;
		memory[16'h6095] <= 8'hca;
		memory[16'h6096] <= 8'h7b;
		memory[16'h6097] <= 8'h36;
		memory[16'h6098] <= 8'h55;
		memory[16'h6099] <= 8'hfb;
		memory[16'h609a] <= 8'h2e;
		memory[16'h609b] <= 8'hea;
		memory[16'h609c] <= 8'h68;
		memory[16'h609d] <= 8'h38;
		memory[16'h609e] <= 8'h13;
		memory[16'h609f] <= 8'h4d;
		memory[16'h60a0] <= 8'h30;
		memory[16'h60a1] <= 8'hc1;
		memory[16'h60a2] <= 8'h40;
		memory[16'h60a3] <= 8'h94;
		memory[16'h60a4] <= 8'h2c;
		memory[16'h60a5] <= 8'h31;
		memory[16'h60a6] <= 8'hc3;
		memory[16'h60a7] <= 8'h3b;
		memory[16'h60a8] <= 8'hfb;
		memory[16'h60a9] <= 8'hbf;
		memory[16'h60aa] <= 8'hb8;
		memory[16'h60ab] <= 8'h77;
		memory[16'h60ac] <= 8'h41;
		memory[16'h60ad] <= 8'he9;
		memory[16'h60ae] <= 8'h45;
		memory[16'h60af] <= 8'h42;
		memory[16'h60b0] <= 8'hef;
		memory[16'h60b1] <= 8'hf;
		memory[16'h60b2] <= 8'h5b;
		memory[16'h60b3] <= 8'hc1;
		memory[16'h60b4] <= 8'hd9;
		memory[16'h60b5] <= 8'hd7;
		memory[16'h60b6] <= 8'hf7;
		memory[16'h60b7] <= 8'h2f;
		memory[16'h60b8] <= 8'hd2;
		memory[16'h60b9] <= 8'h26;
		memory[16'h60ba] <= 8'h19;
		memory[16'h60bb] <= 8'h3b;
		memory[16'h60bc] <= 8'h5e;
		memory[16'h60bd] <= 8'h2c;
		memory[16'h60be] <= 8'h88;
		memory[16'h60bf] <= 8'h8f;
		memory[16'h60c0] <= 8'hed;
		memory[16'h60c1] <= 8'hc8;
		memory[16'h60c2] <= 8'h23;
		memory[16'h60c3] <= 8'h19;
		memory[16'h60c4] <= 8'hfa;
		memory[16'h60c5] <= 8'he6;
		memory[16'h60c6] <= 8'h54;
		memory[16'h60c7] <= 8'hf5;
		memory[16'h60c8] <= 8'ha5;
		memory[16'h60c9] <= 8'hc;
		memory[16'h60ca] <= 8'h6c;
		memory[16'h60cb] <= 8'he6;
		memory[16'h60cc] <= 8'hf6;
		memory[16'h60cd] <= 8'hb1;
		memory[16'h60ce] <= 8'h29;
		memory[16'h60cf] <= 8'he5;
		memory[16'h60d0] <= 8'hc1;
		memory[16'h60d1] <= 8'h84;
		memory[16'h60d2] <= 8'ha7;
		memory[16'h60d3] <= 8'h9a;
		memory[16'h60d4] <= 8'h5b;
		memory[16'h60d5] <= 8'h9e;
		memory[16'h60d6] <= 8'hc9;
		memory[16'h60d7] <= 8'h2e;
		memory[16'h60d8] <= 8'hc4;
		memory[16'h60d9] <= 8'he2;
		memory[16'h60da] <= 8'h69;
		memory[16'h60db] <= 8'h23;
		memory[16'h60dc] <= 8'he;
		memory[16'h60dd] <= 8'hf1;
		memory[16'h60de] <= 8'hb2;
		memory[16'h60df] <= 8'hfb;
		memory[16'h60e0] <= 8'hba;
		memory[16'h60e1] <= 8'hd5;
		memory[16'h60e2] <= 8'h14;
		memory[16'h60e3] <= 8'hb4;
		memory[16'h60e4] <= 8'hbb;
		memory[16'h60e5] <= 8'h69;
		memory[16'h60e6] <= 8'ha9;
		memory[16'h60e7] <= 8'h60;
		memory[16'h60e8] <= 8'h75;
		memory[16'h60e9] <= 8'h16;
		memory[16'h60ea] <= 8'h47;
		memory[16'h60eb] <= 8'h6b;
		memory[16'h60ec] <= 8'hc7;
		memory[16'h60ed] <= 8'h70;
		memory[16'h60ee] <= 8'h51;
		memory[16'h60ef] <= 8'h88;
		memory[16'h60f0] <= 8'hf4;
		memory[16'h60f1] <= 8'hf8;
		memory[16'h60f2] <= 8'h23;
		memory[16'h60f3] <= 8'h50;
		memory[16'h60f4] <= 8'h96;
		memory[16'h60f5] <= 8'hec;
		memory[16'h60f6] <= 8'h7e;
		memory[16'h60f7] <= 8'h5b;
		memory[16'h60f8] <= 8'hcf;
		memory[16'h60f9] <= 8'he7;
		memory[16'h60fa] <= 8'h7e;
		memory[16'h60fb] <= 8'hdd;
		memory[16'h60fc] <= 8'hd8;
		memory[16'h60fd] <= 8'h30;
		memory[16'h60fe] <= 8'hd9;
		memory[16'h60ff] <= 8'h92;
		memory[16'h6100] <= 8'h5;
		memory[16'h6101] <= 8'hed;
		memory[16'h6102] <= 8'h46;
		memory[16'h6103] <= 8'hc0;
		memory[16'h6104] <= 8'h56;
		memory[16'h6105] <= 8'hf0;
		memory[16'h6106] <= 8'h20;
		memory[16'h6107] <= 8'hcc;
		memory[16'h6108] <= 8'h6;
		memory[16'h6109] <= 8'h67;
		memory[16'h610a] <= 8'h37;
		memory[16'h610b] <= 8'hcd;
		memory[16'h610c] <= 8'hd7;
		memory[16'h610d] <= 8'h88;
		memory[16'h610e] <= 8'h56;
		memory[16'h610f] <= 8'hcc;
		memory[16'h6110] <= 8'h80;
		memory[16'h6111] <= 8'h79;
		memory[16'h6112] <= 8'h1c;
		memory[16'h6113] <= 8'h17;
		memory[16'h6114] <= 8'h65;
		memory[16'h6115] <= 8'h9a;
		memory[16'h6116] <= 8'h72;
		memory[16'h6117] <= 8'h34;
		memory[16'h6118] <= 8'h81;
		memory[16'h6119] <= 8'hf0;
		memory[16'h611a] <= 8'h12;
		memory[16'h611b] <= 8'h59;
		memory[16'h611c] <= 8'h20;
		memory[16'h611d] <= 8'heb;
		memory[16'h611e] <= 8'hec;
		memory[16'h611f] <= 8'h25;
		memory[16'h6120] <= 8'hd8;
		memory[16'h6121] <= 8'h32;
		memory[16'h6122] <= 8'he5;
		memory[16'h6123] <= 8'h2f;
		memory[16'h6124] <= 8'h22;
		memory[16'h6125] <= 8'h5;
		memory[16'h6126] <= 8'hfb;
		memory[16'h6127] <= 8'h28;
		memory[16'h6128] <= 8'h6d;
		memory[16'h6129] <= 8'h32;
		memory[16'h612a] <= 8'hf6;
		memory[16'h612b] <= 8'h44;
		memory[16'h612c] <= 8'hbb;
		memory[16'h612d] <= 8'h4c;
		memory[16'h612e] <= 8'h10;
		memory[16'h612f] <= 8'h3b;
		memory[16'h6130] <= 8'hc5;
		memory[16'h6131] <= 8'h2c;
		memory[16'h6132] <= 8'h52;
		memory[16'h6133] <= 8'h2a;
		memory[16'h6134] <= 8'hc6;
		memory[16'h6135] <= 8'hc4;
		memory[16'h6136] <= 8'h5f;
		memory[16'h6137] <= 8'h47;
		memory[16'h6138] <= 8'hb4;
		memory[16'h6139] <= 8'h71;
		memory[16'h613a] <= 8'ha1;
		memory[16'h613b] <= 8'hd4;
		memory[16'h613c] <= 8'h5c;
		memory[16'h613d] <= 8'h8d;
		memory[16'h613e] <= 8'hf9;
		memory[16'h613f] <= 8'h34;
		memory[16'h6140] <= 8'hbf;
		memory[16'h6141] <= 8'hde;
		memory[16'h6142] <= 8'h63;
		memory[16'h6143] <= 8'he2;
		memory[16'h6144] <= 8'he4;
		memory[16'h6145] <= 8'h5e;
		memory[16'h6146] <= 8'ha;
		memory[16'h6147] <= 8'h51;
		memory[16'h6148] <= 8'h91;
		memory[16'h6149] <= 8'h0;
		memory[16'h614a] <= 8'h95;
		memory[16'h614b] <= 8'h4c;
		memory[16'h614c] <= 8'h4c;
		memory[16'h614d] <= 8'ha6;
		memory[16'h614e] <= 8'h87;
		memory[16'h614f] <= 8'h11;
		memory[16'h6150] <= 8'hd2;
		memory[16'h6151] <= 8'hda;
		memory[16'h6152] <= 8'h3c;
		memory[16'h6153] <= 8'h99;
		memory[16'h6154] <= 8'h9e;
		memory[16'h6155] <= 8'h9b;
		memory[16'h6156] <= 8'he0;
		memory[16'h6157] <= 8'h53;
		memory[16'h6158] <= 8'hc;
		memory[16'h6159] <= 8'h81;
		memory[16'h615a] <= 8'h27;
		memory[16'h615b] <= 8'h68;
		memory[16'h615c] <= 8'he;
		memory[16'h615d] <= 8'h21;
		memory[16'h615e] <= 8'h9c;
		memory[16'h615f] <= 8'hce;
		memory[16'h6160] <= 8'hff;
		memory[16'h6161] <= 8'h0;
		memory[16'h6162] <= 8'hb0;
		memory[16'h6163] <= 8'he3;
		memory[16'h6164] <= 8'h5e;
		memory[16'h6165] <= 8'hba;
		memory[16'h6166] <= 8'h34;
		memory[16'h6167] <= 8'hef;
		memory[16'h6168] <= 8'hbb;
		memory[16'h6169] <= 8'hca;
		memory[16'h616a] <= 8'h3b;
		memory[16'h616b] <= 8'h7;
		memory[16'h616c] <= 8'h70;
		memory[16'h616d] <= 8'hc3;
		memory[16'h616e] <= 8'h19;
		memory[16'h616f] <= 8'h42;
		memory[16'h6170] <= 8'h9d;
		memory[16'h6171] <= 8'h55;
		memory[16'h6172] <= 8'hdb;
		memory[16'h6173] <= 8'h3b;
		memory[16'h6174] <= 8'hf0;
		memory[16'h6175] <= 8'hbc;
		memory[16'h6176] <= 8'h8e;
		memory[16'h6177] <= 8'hfc;
		memory[16'h6178] <= 8'h3d;
		memory[16'h6179] <= 8'hb6;
		memory[16'h617a] <= 8'h64;
		memory[16'h617b] <= 8'h4c;
		memory[16'h617c] <= 8'hd7;
		memory[16'h617d] <= 8'h0;
		memory[16'h617e] <= 8'h1a;
		memory[16'h617f] <= 8'hd6;
		memory[16'h6180] <= 8'h0;
		memory[16'h6181] <= 8'hca;
		memory[16'h6182] <= 8'hba;
		memory[16'h6183] <= 8'h5f;
		memory[16'h6184] <= 8'h84;
		memory[16'h6185] <= 8'hee;
		memory[16'h6186] <= 8'h4e;
		memory[16'h6187] <= 8'h3f;
		memory[16'h6188] <= 8'hb8;
		memory[16'h6189] <= 8'h8a;
		memory[16'h618a] <= 8'h47;
		memory[16'h618b] <= 8'h28;
		memory[16'h618c] <= 8'h4d;
		memory[16'h618d] <= 8'h60;
		memory[16'h618e] <= 8'h6b;
		memory[16'h618f] <= 8'hea;
		memory[16'h6190] <= 8'hb5;
		memory[16'h6191] <= 8'h46;
		memory[16'h6192] <= 8'h25;
		memory[16'h6193] <= 8'ha5;
		memory[16'h6194] <= 8'h2;
		memory[16'h6195] <= 8'hb4;
		memory[16'h6196] <= 8'ha1;
		memory[16'h6197] <= 8'h40;
		memory[16'h6198] <= 8'h6a;
		memory[16'h6199] <= 8'h5;
		memory[16'h619a] <= 8'h8c;
		memory[16'h619b] <= 8'h41;
		memory[16'h619c] <= 8'h5;
		memory[16'h619d] <= 8'ha6;
		memory[16'h619e] <= 8'h17;
		memory[16'h619f] <= 8'h6;
		memory[16'h61a0] <= 8'h70;
		memory[16'h61a1] <= 8'hd1;
		memory[16'h61a2] <= 8'h65;
		memory[16'h61a3] <= 8'hf4;
		memory[16'h61a4] <= 8'hc0;
		memory[16'h61a5] <= 8'hb3;
		memory[16'h61a6] <= 8'h34;
		memory[16'h61a7] <= 8'h78;
		memory[16'h61a8] <= 8'h3d;
		memory[16'h61a9] <= 8'h7b;
		memory[16'h61aa] <= 8'ha1;
		memory[16'h61ab] <= 8'h8a;
		memory[16'h61ac] <= 8'hdb;
		memory[16'h61ad] <= 8'hc;
		memory[16'h61ae] <= 8'h74;
		memory[16'h61af] <= 8'h90;
		memory[16'h61b0] <= 8'h52;
		memory[16'h61b1] <= 8'h9a;
		memory[16'h61b2] <= 8'h35;
		memory[16'h61b3] <= 8'h55;
		memory[16'h61b4] <= 8'h4e;
		memory[16'h61b5] <= 8'hd6;
		memory[16'h61b6] <= 8'h95;
		memory[16'h61b7] <= 8'hb8;
		memory[16'h61b8] <= 8'hdb;
		memory[16'h61b9] <= 8'h21;
		memory[16'h61ba] <= 8'hf9;
		memory[16'h61bb] <= 8'he0;
		memory[16'h61bc] <= 8'hc7;
		memory[16'h61bd] <= 8'h10;
		memory[16'h61be] <= 8'he6;
		memory[16'h61bf] <= 8'h37;
		memory[16'h61c0] <= 8'he2;
		memory[16'h61c1] <= 8'h4b;
		memory[16'h61c2] <= 8'h2b;
		memory[16'h61c3] <= 8'ha2;
		memory[16'h61c4] <= 8'hff;
		memory[16'h61c5] <= 8'h5f;
		memory[16'h61c6] <= 8'h1a;
		memory[16'h61c7] <= 8'h3c;
		memory[16'h61c8] <= 8'hda;
		memory[16'h61c9] <= 8'hbb;
		memory[16'h61ca] <= 8'hc7;
		memory[16'h61cb] <= 8'hb5;
		memory[16'h61cc] <= 8'hc7;
		memory[16'h61cd] <= 8'h3b;
		memory[16'h61ce] <= 8'h45;
		memory[16'h61cf] <= 8'h1a;
		memory[16'h61d0] <= 8'hd5;
		memory[16'h61d1] <= 8'h7a;
		memory[16'h61d2] <= 8'h6f;
		memory[16'h61d3] <= 8'h23;
		memory[16'h61d4] <= 8'h50;
		memory[16'h61d5] <= 8'h4;
		memory[16'h61d6] <= 8'hdb;
		memory[16'h61d7] <= 8'h2b;
		memory[16'h61d8] <= 8'h25;
		memory[16'h61d9] <= 8'hd4;
		memory[16'h61da] <= 8'hc;
		memory[16'h61db] <= 8'hec;
		memory[16'h61dc] <= 8'he5;
		memory[16'h61dd] <= 8'hf2;
		memory[16'h61de] <= 8'h23;
		memory[16'h61df] <= 8'hc7;
		memory[16'h61e0] <= 8'h3e;
		memory[16'h61e1] <= 8'h4e;
		memory[16'h61e2] <= 8'h69;
		memory[16'h61e3] <= 8'h3d;
		memory[16'h61e4] <= 8'hae;
		memory[16'h61e5] <= 8'h83;
		memory[16'h61e6] <= 8'h79;
		memory[16'h61e7] <= 8'h88;
		memory[16'h61e8] <= 8'h3f;
		memory[16'h61e9] <= 8'h40;
		memory[16'h61ea] <= 8'h3e;
		memory[16'h61eb] <= 8'h6;
		memory[16'h61ec] <= 8'h7c;
		memory[16'h61ed] <= 8'h83;
		memory[16'h61ee] <= 8'h20;
		memory[16'h61ef] <= 8'h51;
		memory[16'h61f0] <= 8'hfe;
		memory[16'h61f1] <= 8'h8f;
		memory[16'h61f2] <= 8'h75;
		memory[16'h61f3] <= 8'h4e;
		memory[16'h61f4] <= 8'h93;
		memory[16'h61f5] <= 8'h50;
		memory[16'h61f6] <= 8'h7a;
		memory[16'h61f7] <= 8'hb8;
		memory[16'h61f8] <= 8'h25;
		memory[16'h61f9] <= 8'h86;
		memory[16'h61fa] <= 8'ha4;
		memory[16'h61fb] <= 8'ha;
		memory[16'h61fc] <= 8'h78;
		memory[16'h61fd] <= 8'hc7;
		memory[16'h61fe] <= 8'hd1;
		memory[16'h61ff] <= 8'hb6;
		memory[16'h6200] <= 8'h16;
		memory[16'h6201] <= 8'h3a;
		memory[16'h6202] <= 8'hf3;
		memory[16'h6203] <= 8'hc4;
		memory[16'h6204] <= 8'hbd;
		memory[16'h6205] <= 8'h6d;
		memory[16'h6206] <= 8'h4c;
		memory[16'h6207] <= 8'hfc;
		memory[16'h6208] <= 8'had;
		memory[16'h6209] <= 8'h8a;
		memory[16'h620a] <= 8'h3;
		memory[16'h620b] <= 8'h29;
		memory[16'h620c] <= 8'he;
		memory[16'h620d] <= 8'h23;
		memory[16'h620e] <= 8'h7b;
		memory[16'h620f] <= 8'hc;
		memory[16'h6210] <= 8'hb3;
		memory[16'h6211] <= 8'hf0;
		memory[16'h6212] <= 8'h5a;
		memory[16'h6213] <= 8'h46;
		memory[16'h6214] <= 8'h40;
		memory[16'h6215] <= 8'hd4;
		memory[16'h6216] <= 8'hff;
		memory[16'h6217] <= 8'h65;
		memory[16'h6218] <= 8'h5a;
		memory[16'h6219] <= 8'ha3;
		memory[16'h621a] <= 8'h6f;
		memory[16'h621b] <= 8'hd3;
		memory[16'h621c] <= 8'h6b;
		memory[16'h621d] <= 8'h40;
		memory[16'h621e] <= 8'h89;
		memory[16'h621f] <= 8'h81;
		memory[16'h6220] <= 8'h7a;
		memory[16'h6221] <= 8'h7d;
		memory[16'h6222] <= 8'h45;
		memory[16'h6223] <= 8'h38;
		memory[16'h6224] <= 8'hea;
		memory[16'h6225] <= 8'h91;
		memory[16'h6226] <= 8'h34;
		memory[16'h6227] <= 8'h97;
		memory[16'h6228] <= 8'h1c;
		memory[16'h6229] <= 8'h37;
		memory[16'h622a] <= 8'hc1;
		memory[16'h622b] <= 8'h2a;
		memory[16'h622c] <= 8'h5b;
		memory[16'h622d] <= 8'h3c;
		memory[16'h622e] <= 8'h36;
		memory[16'h622f] <= 8'he;
		memory[16'h6230] <= 8'h2c;
		memory[16'h6231] <= 8'h90;
		memory[16'h6232] <= 8'h54;
		memory[16'h6233] <= 8'h6c;
		memory[16'h6234] <= 8'h65;
		memory[16'h6235] <= 8'h53;
		memory[16'h6236] <= 8'hd2;
		memory[16'h6237] <= 8'hbf;
		memory[16'h6238] <= 8'hf7;
		memory[16'h6239] <= 8'h41;
		memory[16'h623a] <= 8'h92;
		memory[16'h623b] <= 8'h62;
		memory[16'h623c] <= 8'h82;
		memory[16'h623d] <= 8'h1c;
		memory[16'h623e] <= 8'he3;
		memory[16'h623f] <= 8'hfc;
		memory[16'h6240] <= 8'h99;
		memory[16'h6241] <= 8'h28;
		memory[16'h6242] <= 8'h34;
		memory[16'h6243] <= 8'h83;
		memory[16'h6244] <= 8'hb9;
		memory[16'h6245] <= 8'h69;
		memory[16'h6246] <= 8'h1a;
		memory[16'h6247] <= 8'hd5;
		memory[16'h6248] <= 8'ha0;
		memory[16'h6249] <= 8'hdb;
		memory[16'h624a] <= 8'hff;
		memory[16'h624b] <= 8'hfb;
		memory[16'h624c] <= 8'h17;
		memory[16'h624d] <= 8'h35;
		memory[16'h624e] <= 8'h9;
		memory[16'h624f] <= 8'h43;
		memory[16'h6250] <= 8'hc6;
		memory[16'h6251] <= 8'h5e;
		memory[16'h6252] <= 8'hb0;
		memory[16'h6253] <= 8'h2b;
		memory[16'h6254] <= 8'hb1;
		memory[16'h6255] <= 8'h82;
		memory[16'h6256] <= 8'hea;
		memory[16'h6257] <= 8'ha8;
		memory[16'h6258] <= 8'hc3;
		memory[16'h6259] <= 8'h7d;
		memory[16'h625a] <= 8'ha;
		memory[16'h625b] <= 8'h45;
		memory[16'h625c] <= 8'h99;
		memory[16'h625d] <= 8'hed;
		memory[16'h625e] <= 8'h42;
		memory[16'h625f] <= 8'h32;
		memory[16'h6260] <= 8'h15;
		memory[16'h6261] <= 8'h76;
		memory[16'h6262] <= 8'hb5;
		memory[16'h6263] <= 8'hcf;
		memory[16'h6264] <= 8'hdf;
		memory[16'h6265] <= 8'hcf;
		memory[16'h6266] <= 8'ha4;
		memory[16'h6267] <= 8'h80;
		memory[16'h6268] <= 8'hab;
		memory[16'h6269] <= 8'ha4;
		memory[16'h626a] <= 8'h7b;
		memory[16'h626b] <= 8'hc2;
		memory[16'h626c] <= 8'hd9;
		memory[16'h626d] <= 8'h85;
		memory[16'h626e] <= 8'h6;
		memory[16'h626f] <= 8'h9f;
		memory[16'h6270] <= 8'he3;
		memory[16'h6271] <= 8'hb6;
		memory[16'h6272] <= 8'hca;
		memory[16'h6273] <= 8'h94;
		memory[16'h6274] <= 8'h38;
		memory[16'h6275] <= 8'hb5;
		memory[16'h6276] <= 8'h3d;
		memory[16'h6277] <= 8'hfb;
		memory[16'h6278] <= 8'h32;
		memory[16'h6279] <= 8'h47;
		memory[16'h627a] <= 8'h41;
		memory[16'h627b] <= 8'hcb;
		memory[16'h627c] <= 8'h35;
		memory[16'h627d] <= 8'h83;
		memory[16'h627e] <= 8'hfd;
		memory[16'h627f] <= 8'h4a;
		memory[16'h6280] <= 8'hf9;
		memory[16'h6281] <= 8'hb2;
		memory[16'h6282] <= 8'h19;
		memory[16'h6283] <= 8'hd9;
		memory[16'h6284] <= 8'h81;
		memory[16'h6285] <= 8'hbe;
		memory[16'h6286] <= 8'h59;
		memory[16'h6287] <= 8'h2c;
		memory[16'h6288] <= 8'h62;
		memory[16'h6289] <= 8'hd4;
		memory[16'h628a] <= 8'hef;
		memory[16'h628b] <= 8'h3b;
		memory[16'h628c] <= 8'h59;
		memory[16'h628d] <= 8'hf5;
		memory[16'h628e] <= 8'hdb;
		memory[16'h628f] <= 8'h3c;
		memory[16'h6290] <= 8'hab;
		memory[16'h6291] <= 8'ha5;
		memory[16'h6292] <= 8'hd1;
		memory[16'h6293] <= 8'he3;
		memory[16'h6294] <= 8'h5a;
		memory[16'h6295] <= 8'he;
		memory[16'h6296] <= 8'hde;
		memory[16'h6297] <= 8'h8c;
		memory[16'h6298] <= 8'h55;
		memory[16'h6299] <= 8'h1f;
		memory[16'h629a] <= 8'h57;
		memory[16'h629b] <= 8'h8a;
		memory[16'h629c] <= 8'ha2;
		memory[16'h629d] <= 8'h54;
		memory[16'h629e] <= 8'hd5;
		memory[16'h629f] <= 8'h9c;
		memory[16'h62a0] <= 8'h6;
		memory[16'h62a1] <= 8'hee;
		memory[16'h62a2] <= 8'h75;
		memory[16'h62a3] <= 8'h88;
		memory[16'h62a4] <= 8'hac;
		memory[16'h62a5] <= 8'hce;
		memory[16'h62a6] <= 8'hb4;
		memory[16'h62a7] <= 8'he;
		memory[16'h62a8] <= 8'ha2;
		memory[16'h62a9] <= 8'ha3;
		memory[16'h62aa] <= 8'h4a;
		memory[16'h62ab] <= 8'hfc;
		memory[16'h62ac] <= 8'h98;
		memory[16'h62ad] <= 8'h25;
		memory[16'h62ae] <= 8'h38;
		memory[16'h62af] <= 8'h43;
		memory[16'h62b0] <= 8'hca;
		memory[16'h62b1] <= 8'h9;
		memory[16'h62b2] <= 8'h26;
		memory[16'h62b3] <= 8'h25;
		memory[16'h62b4] <= 8'h17;
		memory[16'h62b5] <= 8'h5;
		memory[16'h62b6] <= 8'hb1;
		memory[16'h62b7] <= 8'h6d;
		memory[16'h62b8] <= 8'h24;
		memory[16'h62b9] <= 8'h9;
		memory[16'h62ba] <= 8'hf7;
		memory[16'h62bb] <= 8'hc7;
		memory[16'h62bc] <= 8'h5d;
		memory[16'h62bd] <= 8'hcc;
		memory[16'h62be] <= 8'h63;
		memory[16'h62bf] <= 8'h64;
		memory[16'h62c0] <= 8'hbb;
		memory[16'h62c1] <= 8'hd8;
		memory[16'h62c2] <= 8'hec;
		memory[16'h62c3] <= 8'h67;
		memory[16'h62c4] <= 8'ha6;
		memory[16'h62c5] <= 8'ha0;
		memory[16'h62c6] <= 8'h76;
		memory[16'h62c7] <= 8'h48;
		memory[16'h62c8] <= 8'h44;
		memory[16'h62c9] <= 8'hc0;
		memory[16'h62ca] <= 8'h44;
		memory[16'h62cb] <= 8'hdc;
		memory[16'h62cc] <= 8'he5;
		memory[16'h62cd] <= 8'h7d;
		memory[16'h62ce] <= 8'h20;
		memory[16'h62cf] <= 8'haf;
		memory[16'h62d0] <= 8'h86;
		memory[16'h62d1] <= 8'h46;
		memory[16'h62d2] <= 8'hd4;
		memory[16'h62d3] <= 8'h9e;
		memory[16'h62d4] <= 8'h4b;
		memory[16'h62d5] <= 8'h86;
		memory[16'h62d6] <= 8'hb;
		memory[16'h62d7] <= 8'h70;
		memory[16'h62d8] <= 8'h8f;
		memory[16'h62d9] <= 8'h2;
		memory[16'h62da] <= 8'h37;
		memory[16'h62db] <= 8'hec;
		memory[16'h62dc] <= 8'hcf;
		memory[16'h62dd] <= 8'h9a;
		memory[16'h62de] <= 8'h50;
		memory[16'h62df] <= 8'h8a;
		memory[16'h62e0] <= 8'h72;
		memory[16'h62e1] <= 8'h3c;
		memory[16'h62e2] <= 8'hf1;
		memory[16'h62e3] <= 8'h18;
		memory[16'h62e4] <= 8'hdd;
		memory[16'h62e5] <= 8'h67;
		memory[16'h62e6] <= 8'h60;
		memory[16'h62e7] <= 8'h21;
		memory[16'h62e8] <= 8'h27;
		memory[16'h62e9] <= 8'ha5;
		memory[16'h62ea] <= 8'hfd;
		memory[16'h62eb] <= 8'hc;
		memory[16'h62ec] <= 8'h22;
		memory[16'h62ed] <= 8'h1d;
		memory[16'h62ee] <= 8'hbc;
		memory[16'h62ef] <= 8'ha8;
		memory[16'h62f0] <= 8'h64;
		memory[16'h62f1] <= 8'h90;
		memory[16'h62f2] <= 8'h46;
		memory[16'h62f3] <= 8'haf;
		memory[16'h62f4] <= 8'h16;
		memory[16'h62f5] <= 8'h51;
		memory[16'h62f6] <= 8'h1f;
		memory[16'h62f7] <= 8'ha5;
		memory[16'h62f8] <= 8'h54;
		memory[16'h62f9] <= 8'h56;
		memory[16'h62fa] <= 8'h92;
		memory[16'h62fb] <= 8'h23;
		memory[16'h62fc] <= 8'hf0;
		memory[16'h62fd] <= 8'he2;
		memory[16'h62fe] <= 8'had;
		memory[16'h62ff] <= 8'h62;
		memory[16'h6300] <= 8'h1f;
		memory[16'h6301] <= 8'h9e;
		memory[16'h6302] <= 8'h7a;
		memory[16'h6303] <= 8'hfc;
		memory[16'h6304] <= 8'h6;
		memory[16'h6305] <= 8'hdb;
		memory[16'h6306] <= 8'h1d;
		memory[16'h6307] <= 8'h2d;
		memory[16'h6308] <= 8'h80;
		memory[16'h6309] <= 8'h1a;
		memory[16'h630a] <= 8'h3a;
		memory[16'h630b] <= 8'ha2;
		memory[16'h630c] <= 8'h38;
		memory[16'h630d] <= 8'hf6;
		memory[16'h630e] <= 8'h4a;
		memory[16'h630f] <= 8'h9c;
		memory[16'h6310] <= 8'h86;
		memory[16'h6311] <= 8'h91;
		memory[16'h6312] <= 8'h4b;
		memory[16'h6313] <= 8'h9d;
		memory[16'h6314] <= 8'he2;
		memory[16'h6315] <= 8'h6b;
		memory[16'h6316] <= 8'h42;
		memory[16'h6317] <= 8'h36;
		memory[16'h6318] <= 8'hc1;
		memory[16'h6319] <= 8'hd4;
		memory[16'h631a] <= 8'h59;
		memory[16'h631b] <= 8'hb2;
		memory[16'h631c] <= 8'hb7;
		memory[16'h631d] <= 8'h6;
		memory[16'h631e] <= 8'h14;
		memory[16'h631f] <= 8'hd6;
		memory[16'h6320] <= 8'ha5;
		memory[16'h6321] <= 8'h8f;
		memory[16'h6322] <= 8'hd2;
		memory[16'h6323] <= 8'hab;
		memory[16'h6324] <= 8'h6a;
		memory[16'h6325] <= 8'hef;
		memory[16'h6326] <= 8'hd8;
		memory[16'h6327] <= 8'hea;
		memory[16'h6328] <= 8'h9;
		memory[16'h6329] <= 8'h12;
		memory[16'h632a] <= 8'h8c;
		memory[16'h632b] <= 8'h41;
		memory[16'h632c] <= 8'h8;
		memory[16'h632d] <= 8'hd6;
		memory[16'h632e] <= 8'hdd;
		memory[16'h632f] <= 8'h8f;
		memory[16'h6330] <= 8'h67;
		memory[16'h6331] <= 8'h29;
		memory[16'h6332] <= 8'h2c;
		memory[16'h6333] <= 8'h4a;
		memory[16'h6334] <= 8'h94;
		memory[16'h6335] <= 8'h6e;
		memory[16'h6336] <= 8'h80;
		memory[16'h6337] <= 8'h55;
		memory[16'h6338] <= 8'h43;
		memory[16'h6339] <= 8'hda;
		memory[16'h633a] <= 8'h7;
		memory[16'h633b] <= 8'hfa;
		memory[16'h633c] <= 8'he0;
		memory[16'h633d] <= 8'h1c;
		memory[16'h633e] <= 8'hd0;
		memory[16'h633f] <= 8'h85;
		memory[16'h6340] <= 8'hab;
		memory[16'h6341] <= 8'ha2;
		memory[16'h6342] <= 8'h30;
		memory[16'h6343] <= 8'h15;
		memory[16'h6344] <= 8'h91;
		memory[16'h6345] <= 8'h9;
		memory[16'h6346] <= 8'hff;
		memory[16'h6347] <= 8'h9a;
		memory[16'h6348] <= 8'h1b;
		memory[16'h6349] <= 8'h8b;
		memory[16'h634a] <= 8'hdc;
		memory[16'h634b] <= 8'h24;
		memory[16'h634c] <= 8'h61;
		memory[16'h634d] <= 8'hb9;
		memory[16'h634e] <= 8'hb3;
		memory[16'h634f] <= 8'hc9;
		memory[16'h6350] <= 8'he2;
		memory[16'h6351] <= 8'hdf;
		memory[16'h6352] <= 8'h13;
		memory[16'h6353] <= 8'h76;
		memory[16'h6354] <= 8'h4d;
		memory[16'h6355] <= 8'h93;
		memory[16'h6356] <= 8'hcc;
		memory[16'h6357] <= 8'h90;
		memory[16'h6358] <= 8'h6d;
		memory[16'h6359] <= 8'hd3;
		memory[16'h635a] <= 8'h8a;
		memory[16'h635b] <= 8'h4e;
		memory[16'h635c] <= 8'hef;
		memory[16'h635d] <= 8'h5a;
		memory[16'h635e] <= 8'hd3;
		memory[16'h635f] <= 8'h9a;
		memory[16'h6360] <= 8'hfc;
		memory[16'h6361] <= 8'h4;
		memory[16'h6362] <= 8'haf;
		memory[16'h6363] <= 8'h8d;
		memory[16'h6364] <= 8'hd;
		memory[16'h6365] <= 8'hae;
		memory[16'h6366] <= 8'h28;
		memory[16'h6367] <= 8'h28;
		memory[16'h6368] <= 8'h39;
		memory[16'h6369] <= 8'h4;
		memory[16'h636a] <= 8'h4c;
		memory[16'h636b] <= 8'h9b;
		memory[16'h636c] <= 8'hbd;
		memory[16'h636d] <= 8'hff;
		memory[16'h636e] <= 8'h64;
		memory[16'h636f] <= 8'ha0;
		memory[16'h6370] <= 8'hde;
		memory[16'h6371] <= 8'h77;
		memory[16'h6372] <= 8'h16;
		memory[16'h6373] <= 8'h2c;
		memory[16'h6374] <= 8'ha;
		memory[16'h6375] <= 8'he2;
		memory[16'h6376] <= 8'hbc;
		memory[16'h6377] <= 8'h78;
		memory[16'h6378] <= 8'hb6;
		memory[16'h6379] <= 8'h47;
		memory[16'h637a] <= 8'hc6;
		memory[16'h637b] <= 8'ha5;
		memory[16'h637c] <= 8'ha1;
		memory[16'h637d] <= 8'h99;
		memory[16'h637e] <= 8'h40;
		memory[16'h637f] <= 8'h9e;
		memory[16'h6380] <= 8'h9d;
		memory[16'h6381] <= 8'hef;
		memory[16'h6382] <= 8'h2b;
		memory[16'h6383] <= 8'haa;
		memory[16'h6384] <= 8'h9e;
		memory[16'h6385] <= 8'h53;
		memory[16'h6386] <= 8'hd3;
		memory[16'h6387] <= 8'hd7;
		memory[16'h6388] <= 8'h57;
		memory[16'h6389] <= 8'h1f;
		memory[16'h638a] <= 8'h72;
		memory[16'h638b] <= 8'h15;
		memory[16'h638c] <= 8'h1f;
		memory[16'h638d] <= 8'hd6;
		memory[16'h638e] <= 8'hb5;
		memory[16'h638f] <= 8'hfd;
		memory[16'h6390] <= 8'h4d;
		memory[16'h6391] <= 8'hcb;
		memory[16'h6392] <= 8'h29;
		memory[16'h6393] <= 8'h58;
		memory[16'h6394] <= 8'hae;
		memory[16'h6395] <= 8'he6;
		memory[16'h6396] <= 8'hd0;
		memory[16'h6397] <= 8'h64;
		memory[16'h6398] <= 8'h2d;
		memory[16'h6399] <= 8'h96;
		memory[16'h639a] <= 8'h9;
		memory[16'h639b] <= 8'hce;
		memory[16'h639c] <= 8'h2f;
		memory[16'h639d] <= 8'h49;
		memory[16'h639e] <= 8'h6c;
		memory[16'h639f] <= 8'hcd;
		memory[16'h63a0] <= 8'h39;
		memory[16'h63a1] <= 8'h98;
		memory[16'h63a2] <= 8'h77;
		memory[16'h63a3] <= 8'hd7;
		memory[16'h63a4] <= 8'heb;
		memory[16'h63a5] <= 8'h4a;
		memory[16'h63a6] <= 8'hae;
		memory[16'h63a7] <= 8'h43;
		memory[16'h63a8] <= 8'h6a;
		memory[16'h63a9] <= 8'h21;
		memory[16'h63aa] <= 8'h58;
		memory[16'h63ab] <= 8'h89;
		memory[16'h63ac] <= 8'hf7;
		memory[16'h63ad] <= 8'hd;
		memory[16'h63ae] <= 8'h86;
		memory[16'h63af] <= 8'h45;
		memory[16'h63b0] <= 8'hd8;
		memory[16'h63b1] <= 8'hb0;
		memory[16'h63b2] <= 8'h9d;
		memory[16'h63b3] <= 8'h86;
		memory[16'h63b4] <= 8'h96;
		memory[16'h63b5] <= 8'h6d;
		memory[16'h63b6] <= 8'hea;
		memory[16'h63b7] <= 8'hc3;
		memory[16'h63b8] <= 8'h3;
		memory[16'h63b9] <= 8'hf4;
		memory[16'h63ba] <= 8'h91;
		memory[16'h63bb] <= 8'h32;
		memory[16'h63bc] <= 8'h3d;
		memory[16'h63bd] <= 8'hfe;
		memory[16'h63be] <= 8'hff;
		memory[16'h63bf] <= 8'h76;
		memory[16'h63c0] <= 8'h96;
		memory[16'h63c1] <= 8'h77;
		memory[16'h63c2] <= 8'h4d;
		memory[16'h63c3] <= 8'h81;
		memory[16'h63c4] <= 8'hc1;
		memory[16'h63c5] <= 8'hfc;
		memory[16'h63c6] <= 8'hc4;
		memory[16'h63c7] <= 8'h2b;
		memory[16'h63c8] <= 8'h1d;
		memory[16'h63c9] <= 8'h1c;
		memory[16'h63ca] <= 8'hb4;
		memory[16'h63cb] <= 8'h14;
		memory[16'h63cc] <= 8'h29;
		memory[16'h63cd] <= 8'h3b;
		memory[16'h63ce] <= 8'h59;
		memory[16'h63cf] <= 8'h2;
		memory[16'h63d0] <= 8'heb;
		memory[16'h63d1] <= 8'hf6;
		memory[16'h63d2] <= 8'h88;
		memory[16'h63d3] <= 8'h81;
		memory[16'h63d4] <= 8'h63;
		memory[16'h63d5] <= 8'h73;
		memory[16'h63d6] <= 8'h44;
		memory[16'h63d7] <= 8'h66;
		memory[16'h63d8] <= 8'h67;
		memory[16'h63d9] <= 8'hd5;
		memory[16'h63da] <= 8'h99;
		memory[16'h63db] <= 8'ha4;
		memory[16'h63dc] <= 8'hd3;
		memory[16'h63dd] <= 8'h98;
		memory[16'h63de] <= 8'h1b;
		memory[16'h63df] <= 8'h69;
		memory[16'h63e0] <= 8'hf;
		memory[16'h63e1] <= 8'h68;
		memory[16'h63e2] <= 8'heb;
		memory[16'h63e3] <= 8'hd1;
		memory[16'h63e4] <= 8'h64;
		memory[16'h63e5] <= 8'haf;
		memory[16'h63e6] <= 8'hfc;
		memory[16'h63e7] <= 8'h81;
		memory[16'h63e8] <= 8'hcc;
		memory[16'h63e9] <= 8'hb1;
		memory[16'h63ea] <= 8'h96;
		memory[16'h63eb] <= 8'hf5;
		memory[16'h63ec] <= 8'hec;
		memory[16'h63ed] <= 8'hef;
		memory[16'h63ee] <= 8'hf7;
		memory[16'h63ef] <= 8'hd7;
		memory[16'h63f0] <= 8'he6;
		memory[16'h63f1] <= 8'h80;
		memory[16'h63f2] <= 8'h58;
		memory[16'h63f3] <= 8'h49;
		memory[16'h63f4] <= 8'hf3;
		memory[16'h63f5] <= 8'h9c;
		memory[16'h63f6] <= 8'hb0;
		memory[16'h63f7] <= 8'h5a;
		memory[16'h63f8] <= 8'h71;
		memory[16'h63f9] <= 8'h49;
		memory[16'h63fa] <= 8'hfe;
		memory[16'h63fb] <= 8'h45;
		memory[16'h63fc] <= 8'he1;
		memory[16'h63fd] <= 8'h19;
		memory[16'h63fe] <= 8'hae;
		memory[16'h63ff] <= 8'hf1;
		memory[16'h6400] <= 8'h82;
		memory[16'h6401] <= 8'h99;
		memory[16'h6402] <= 8'hc2;
		memory[16'h6403] <= 8'he6;
		memory[16'h6404] <= 8'h49;
		memory[16'h6405] <= 8'hbe;
		memory[16'h6406] <= 8'h68;
		memory[16'h6407] <= 8'h15;
		memory[16'h6408] <= 8'h6f;
		memory[16'h6409] <= 8'hfe;
		memory[16'h640a] <= 8'ha;
		memory[16'h640b] <= 8'h5b;
		memory[16'h640c] <= 8'hed;
		memory[16'h640d] <= 8'h2;
		memory[16'h640e] <= 8'h32;
		memory[16'h640f] <= 8'hd3;
		memory[16'h6410] <= 8'h82;
		memory[16'h6411] <= 8'h8a;
		memory[16'h6412] <= 8'h1d;
		memory[16'h6413] <= 8'h75;
		memory[16'h6414] <= 8'h26;
		memory[16'h6415] <= 8'hcd;
		memory[16'h6416] <= 8'hcf;
		memory[16'h6417] <= 8'h98;
		memory[16'h6418] <= 8'h16;
		memory[16'h6419] <= 8'hcd;
		memory[16'h641a] <= 8'hdd;
		memory[16'h641b] <= 8'hf7;
		memory[16'h641c] <= 8'he7;
		memory[16'h641d] <= 8'h8b;
		memory[16'h641e] <= 8'he8;
		memory[16'h641f] <= 8'h69;
		memory[16'h6420] <= 8'h25;
		memory[16'h6421] <= 8'haa;
		memory[16'h6422] <= 8'h4f;
		memory[16'h6423] <= 8'h6e;
		memory[16'h6424] <= 8'h69;
		memory[16'h6425] <= 8'hb7;
		memory[16'h6426] <= 8'h83;
		memory[16'h6427] <= 8'hd8;
		memory[16'h6428] <= 8'hb5;
		memory[16'h6429] <= 8'h8d;
		memory[16'h642a] <= 8'h34;
		memory[16'h642b] <= 8'ha3;
		memory[16'h642c] <= 8'h8f;
		memory[16'h642d] <= 8'h66;
		memory[16'h642e] <= 8'h76;
		memory[16'h642f] <= 8'h11;
		memory[16'h6430] <= 8'hf1;
		memory[16'h6431] <= 8'h93;
		memory[16'h6432] <= 8'h86;
		memory[16'h6433] <= 8'h17;
		memory[16'h6434] <= 8'h60;
		memory[16'h6435] <= 8'h55;
		memory[16'h6436] <= 8'haf;
		memory[16'h6437] <= 8'h76;
		memory[16'h6438] <= 8'h23;
		memory[16'h6439] <= 8'h8c;
		memory[16'h643a] <= 8'h6e;
		memory[16'h643b] <= 8'ha;
		memory[16'h643c] <= 8'h18;
		memory[16'h643d] <= 8'h56;
		memory[16'h643e] <= 8'h73;
		memory[16'h643f] <= 8'h3d;
		memory[16'h6440] <= 8'h1;
		memory[16'h6441] <= 8'hc2;
		memory[16'h6442] <= 8'hab;
		memory[16'h6443] <= 8'h6a;
		memory[16'h6444] <= 8'h7a;
		memory[16'h6445] <= 8'h2e;
		memory[16'h6446] <= 8'h42;
		memory[16'h6447] <= 8'h2f;
		memory[16'h6448] <= 8'hbb;
		memory[16'h6449] <= 8'h76;
		memory[16'h644a] <= 8'hd2;
		memory[16'h644b] <= 8'h4b;
		memory[16'h644c] <= 8'hdd;
		memory[16'h644d] <= 8'h49;
		memory[16'h644e] <= 8'h5c;
		memory[16'h644f] <= 8'hce;
		memory[16'h6450] <= 8'hdc;
		memory[16'h6451] <= 8'he3;
		memory[16'h6452] <= 8'he5;
		memory[16'h6453] <= 8'h3d;
		memory[16'h6454] <= 8'h38;
		memory[16'h6455] <= 8'h95;
		memory[16'h6456] <= 8'hb3;
		memory[16'h6457] <= 8'h5b;
		memory[16'h6458] <= 8'h21;
		memory[16'h6459] <= 8'h21;
		memory[16'h645a] <= 8'h65;
		memory[16'h645b] <= 8'h39;
		memory[16'h645c] <= 8'h78;
		memory[16'h645d] <= 8'hd8;
		memory[16'h645e] <= 8'h76;
		memory[16'h645f] <= 8'h79;
		memory[16'h6460] <= 8'h9b;
		memory[16'h6461] <= 8'h21;
		memory[16'h6462] <= 8'he3;
		memory[16'h6463] <= 8'h15;
		memory[16'h6464] <= 8'h4f;
		memory[16'h6465] <= 8'h25;
		memory[16'h6466] <= 8'h44;
		memory[16'h6467] <= 8'hb;
		memory[16'h6468] <= 8'h9c;
		memory[16'h6469] <= 8'h17;
		memory[16'h646a] <= 8'h56;
		memory[16'h646b] <= 8'h79;
		memory[16'h646c] <= 8'h60;
		memory[16'h646d] <= 8'hb2;
		memory[16'h646e] <= 8'h47;
		memory[16'h646f] <= 8'h3c;
		memory[16'h6470] <= 8'h95;
		memory[16'h6471] <= 8'h2c;
		memory[16'h6472] <= 8'h79;
		memory[16'h6473] <= 8'hce;
		memory[16'h6474] <= 8'hc1;
		memory[16'h6475] <= 8'h2d;
		memory[16'h6476] <= 8'h29;
		memory[16'h6477] <= 8'he3;
		memory[16'h6478] <= 8'h4e;
		memory[16'h6479] <= 8'h8f;
		memory[16'h647a] <= 8'h1c;
		memory[16'h647b] <= 8'hc6;
		memory[16'h647c] <= 8'h67;
		memory[16'h647d] <= 8'h93;
		memory[16'h647e] <= 8'h3f;
		memory[16'h647f] <= 8'h2;
		memory[16'h6480] <= 8'hb4;
		memory[16'h6481] <= 8'h22;
		memory[16'h6482] <= 8'h17;
		memory[16'h6483] <= 8'h4;
		memory[16'h6484] <= 8'h48;
		memory[16'h6485] <= 8'h5c;
		memory[16'h6486] <= 8'hf;
		memory[16'h6487] <= 8'he4;
		memory[16'h6488] <= 8'h73;
		memory[16'h6489] <= 8'h65;
		memory[16'h648a] <= 8'h5d;
		memory[16'h648b] <= 8'hd3;
		memory[16'h648c] <= 8'h17;
		memory[16'h648d] <= 8'ha4;
		memory[16'h648e] <= 8'hf;
		memory[16'h648f] <= 8'had;
		memory[16'h6490] <= 8'hd0;
		memory[16'h6491] <= 8'h89;
		memory[16'h6492] <= 8'h7b;
		memory[16'h6493] <= 8'h92;
		memory[16'h6494] <= 8'hb6;
		memory[16'h6495] <= 8'ha4;
		memory[16'h6496] <= 8'h75;
		memory[16'h6497] <= 8'h4;
		memory[16'h6498] <= 8'h33;
		memory[16'h6499] <= 8'h91;
		memory[16'h649a] <= 8'hcb;
		memory[16'h649b] <= 8'h9b;
		memory[16'h649c] <= 8'h24;
		memory[16'h649d] <= 8'ha;
		memory[16'h649e] <= 8'h9d;
		memory[16'h649f] <= 8'hd9;
		memory[16'h64a0] <= 8'h2d;
		memory[16'h64a1] <= 8'hb5;
		memory[16'h64a2] <= 8'hdd;
		memory[16'h64a3] <= 8'h75;
		memory[16'h64a4] <= 8'h11;
		memory[16'h64a5] <= 8'hec;
		memory[16'h64a6] <= 8'h59;
		memory[16'h64a7] <= 8'h84;
		memory[16'h64a8] <= 8'h51;
		memory[16'h64a9] <= 8'hb6;
		memory[16'h64aa] <= 8'h57;
		memory[16'h64ab] <= 8'h68;
		memory[16'h64ac] <= 8'h5a;
		memory[16'h64ad] <= 8'h66;
		memory[16'h64ae] <= 8'h15;
		memory[16'h64af] <= 8'h2a;
		memory[16'h64b0] <= 8'hef;
		memory[16'h64b1] <= 8'h90;
		memory[16'h64b2] <= 8'hbc;
		memory[16'h64b3] <= 8'ha5;
		memory[16'h64b4] <= 8'h35;
		memory[16'h64b5] <= 8'h31;
		memory[16'h64b6] <= 8'haa;
		memory[16'h64b7] <= 8'h68;
		memory[16'h64b8] <= 8'hc3;
		memory[16'h64b9] <= 8'h75;
		memory[16'h64ba] <= 8'h3;
		memory[16'h64bb] <= 8'he7;
		memory[16'h64bc] <= 8'h7f;
		memory[16'h64bd] <= 8'ha1;
		memory[16'h64be] <= 8'hc0;
		memory[16'h64bf] <= 8'hac;
		memory[16'h64c0] <= 8'h56;
		memory[16'h64c1] <= 8'h9d;
		memory[16'h64c2] <= 8'h21;
		memory[16'h64c3] <= 8'h67;
		memory[16'h64c4] <= 8'h89;
		memory[16'h64c5] <= 8'h7a;
		memory[16'h64c6] <= 8'heb;
		memory[16'h64c7] <= 8'hda;
		memory[16'h64c8] <= 8'h30;
		memory[16'h64c9] <= 8'h42;
		memory[16'h64ca] <= 8'h43;
		memory[16'h64cb] <= 8'h8a;
		memory[16'h64cc] <= 8'ha8;
		memory[16'h64cd] <= 8'h58;
		memory[16'h64ce] <= 8'hb5;
		memory[16'h64cf] <= 8'h98;
		memory[16'h64d0] <= 8'he9;
		memory[16'h64d1] <= 8'h71;
		memory[16'h64d2] <= 8'h3d;
		memory[16'h64d3] <= 8'h1e;
		memory[16'h64d4] <= 8'ha3;
		memory[16'h64d5] <= 8'he7;
		memory[16'h64d6] <= 8'h86;
		memory[16'h64d7] <= 8'h66;
		memory[16'h64d8] <= 8'h5c;
		memory[16'h64d9] <= 8'h8a;
		memory[16'h64da] <= 8'h4d;
		memory[16'h64db] <= 8'hdc;
		memory[16'h64dc] <= 8'h2b;
		memory[16'h64dd] <= 8'he;
		memory[16'h64de] <= 8'h88;
		memory[16'h64df] <= 8'h81;
		memory[16'h64e0] <= 8'hab;
		memory[16'h64e1] <= 8'haa;
		memory[16'h64e2] <= 8'he8;
		memory[16'h64e3] <= 8'h35;
		memory[16'h64e4] <= 8'h24;
		memory[16'h64e5] <= 8'hd3;
		memory[16'h64e6] <= 8'hf;
		memory[16'h64e7] <= 8'h55;
		memory[16'h64e8] <= 8'h15;
		memory[16'h64e9] <= 8'h52;
		memory[16'h64ea] <= 8'hdf;
		memory[16'h64eb] <= 8'hbd;
		memory[16'h64ec] <= 8'hab;
		memory[16'h64ed] <= 8'h94;
		memory[16'h64ee] <= 8'h55;
		memory[16'h64ef] <= 8'h94;
		memory[16'h64f0] <= 8'h6;
		memory[16'h64f1] <= 8'h93;
		memory[16'h64f2] <= 8'hb2;
		memory[16'h64f3] <= 8'ha9;
		memory[16'h64f4] <= 8'h7a;
		memory[16'h64f5] <= 8'h38;
		memory[16'h64f6] <= 8'hf;
		memory[16'h64f7] <= 8'hd7;
		memory[16'h64f8] <= 8'hc2;
		memory[16'h64f9] <= 8'h5c;
		memory[16'h64fa] <= 8'hb3;
		memory[16'h64fb] <= 8'hed;
		memory[16'h64fc] <= 8'h6a;
		memory[16'h64fd] <= 8'h3b;
		memory[16'h64fe] <= 8'h6e;
		memory[16'h64ff] <= 8'h16;
		memory[16'h6500] <= 8'he5;
		memory[16'h6501] <= 8'h56;
		memory[16'h6502] <= 8'h4b;
		memory[16'h6503] <= 8'ha;
		memory[16'h6504] <= 8'h29;
		memory[16'h6505] <= 8'h5a;
		memory[16'h6506] <= 8'h5f;
		memory[16'h6507] <= 8'h3e;
		memory[16'h6508] <= 8'had;
		memory[16'h6509] <= 8'h3e;
		memory[16'h650a] <= 8'hfc;
		memory[16'h650b] <= 8'h58;
		memory[16'h650c] <= 8'hd3;
		memory[16'h650d] <= 8'h51;
		memory[16'h650e] <= 8'hec;
		memory[16'h650f] <= 8'hd9;
		memory[16'h6510] <= 8'he4;
		memory[16'h6511] <= 8'h9e;
		memory[16'h6512] <= 8'h82;
		memory[16'h6513] <= 8'h5f;
		memory[16'h6514] <= 8'hd6;
		memory[16'h6515] <= 8'h91;
		memory[16'h6516] <= 8'h36;
		memory[16'h6517] <= 8'h99;
		memory[16'h6518] <= 8'hed;
		memory[16'h6519] <= 8'he9;
		memory[16'h651a] <= 8'h86;
		memory[16'h651b] <= 8'h58;
		memory[16'h651c] <= 8'h24;
		memory[16'h651d] <= 8'hf5;
		memory[16'h651e] <= 8'h6e;
		memory[16'h651f] <= 8'ha;
		memory[16'h6520] <= 8'h4b;
		memory[16'h6521] <= 8'hb9;
		memory[16'h6522] <= 8'h14;
		memory[16'h6523] <= 8'h75;
		memory[16'h6524] <= 8'h13;
		memory[16'h6525] <= 8'h73;
		memory[16'h6526] <= 8'hb3;
		memory[16'h6527] <= 8'hc0;
		memory[16'h6528] <= 8'hb1;
		memory[16'h6529] <= 8'haf;
		memory[16'h652a] <= 8'h18;
		memory[16'h652b] <= 8'h84;
		memory[16'h652c] <= 8'h1;
		memory[16'h652d] <= 8'h4;
		memory[16'h652e] <= 8'h5d;
		memory[16'h652f] <= 8'he5;
		memory[16'h6530] <= 8'ha2;
		memory[16'h6531] <= 8'hdf;
		memory[16'h6532] <= 8'h44;
		memory[16'h6533] <= 8'h79;
		memory[16'h6534] <= 8'h70;
		memory[16'h6535] <= 8'h7a;
		memory[16'h6536] <= 8'h12;
		memory[16'h6537] <= 8'h5e;
		memory[16'h6538] <= 8'h63;
		memory[16'h6539] <= 8'h98;
		memory[16'h653a] <= 8'hb6;
		memory[16'h653b] <= 8'h88;
		memory[16'h653c] <= 8'h8d;
		memory[16'h653d] <= 8'h24;
		memory[16'h653e] <= 8'h92;
		memory[16'h653f] <= 8'hd9;
		memory[16'h6540] <= 8'hdd;
		memory[16'h6541] <= 8'ha6;
		memory[16'h6542] <= 8'h4e;
		memory[16'h6543] <= 8'hf0;
		memory[16'h6544] <= 8'h19;
		memory[16'h6545] <= 8'h1;
		memory[16'h6546] <= 8'hb1;
		memory[16'h6547] <= 8'hca;
		memory[16'h6548] <= 8'hb1;
		memory[16'h6549] <= 8'hc9;
		memory[16'h654a] <= 8'h4f;
		memory[16'h654b] <= 8'hb2;
		memory[16'h654c] <= 8'hce;
		memory[16'h654d] <= 8'hac;
		memory[16'h654e] <= 8'h97;
		memory[16'h654f] <= 8'h70;
		memory[16'h6550] <= 8'h8c;
		memory[16'h6551] <= 8'hdc;
		memory[16'h6552] <= 8'he9;
		memory[16'h6553] <= 8'hfc;
		memory[16'h6554] <= 8'h56;
		memory[16'h6555] <= 8'hfb;
		memory[16'h6556] <= 8'h5a;
		memory[16'h6557] <= 8'hba;
		memory[16'h6558] <= 8'h94;
		memory[16'h6559] <= 8'h10;
		memory[16'h655a] <= 8'h42;
		memory[16'h655b] <= 8'h21;
		memory[16'h655c] <= 8'h34;
		memory[16'h655d] <= 8'hd4;
		memory[16'h655e] <= 8'hfa;
		memory[16'h655f] <= 8'h11;
		memory[16'h6560] <= 8'h7a;
		memory[16'h6561] <= 8'h48;
		memory[16'h6562] <= 8'h2;
		memory[16'h6563] <= 8'h93;
		memory[16'h6564] <= 8'h4a;
		memory[16'h6565] <= 8'hb3;
		memory[16'h6566] <= 8'h5d;
		memory[16'h6567] <= 8'hfb;
		memory[16'h6568] <= 8'h7c;
		memory[16'h6569] <= 8'hac;
		memory[16'h656a] <= 8'had;
		memory[16'h656b] <= 8'h4a;
		memory[16'h656c] <= 8'h59;
		memory[16'h656d] <= 8'h44;
		memory[16'h656e] <= 8'hbb;
		memory[16'h656f] <= 8'he5;
		memory[16'h6570] <= 8'h20;
		memory[16'h6571] <= 8'ha4;
		memory[16'h6572] <= 8'he1;
		memory[16'h6573] <= 8'h77;
		memory[16'h6574] <= 8'ha0;
		memory[16'h6575] <= 8'h3c;
		memory[16'h6576] <= 8'h31;
		memory[16'h6577] <= 8'h34;
		memory[16'h6578] <= 8'h4c;
		memory[16'h6579] <= 8'h73;
		memory[16'h657a] <= 8'h55;
		memory[16'h657b] <= 8'h81;
		memory[16'h657c] <= 8'h47;
		memory[16'h657d] <= 8'h50;
		memory[16'h657e] <= 8'h92;
		memory[16'h657f] <= 8'hc1;
		memory[16'h6580] <= 8'h98;
		memory[16'h6581] <= 8'h94;
		memory[16'h6582] <= 8'h54;
		memory[16'h6583] <= 8'he2;
		memory[16'h6584] <= 8'h47;
		memory[16'h6585] <= 8'hb1;
		memory[16'h6586] <= 8'hdd;
		memory[16'h6587] <= 8'hc4;
		memory[16'h6588] <= 8'h5e;
		memory[16'h6589] <= 8'h8a;
		memory[16'h658a] <= 8'he;
		memory[16'h658b] <= 8'hb7;
		memory[16'h658c] <= 8'hcf;
		memory[16'h658d] <= 8'hc9;
		memory[16'h658e] <= 8'h9c;
		memory[16'h658f] <= 8'hef;
		memory[16'h6590] <= 8'h6e;
		memory[16'h6591] <= 8'h7d;
		memory[16'h6592] <= 8'h66;
		memory[16'h6593] <= 8'he;
		memory[16'h6594] <= 8'hb9;
		memory[16'h6595] <= 8'h97;
		memory[16'h6596] <= 8'h42;
		memory[16'h6597] <= 8'h6;
		memory[16'h6598] <= 8'ha;
		memory[16'h6599] <= 8'h97;
		memory[16'h659a] <= 8'h87;
		memory[16'h659b] <= 8'h51;
		memory[16'h659c] <= 8'he7;
		memory[16'h659d] <= 8'h19;
		memory[16'h659e] <= 8'h12;
		memory[16'h659f] <= 8'h80;
		memory[16'h65a0] <= 8'hae;
		memory[16'h65a1] <= 8'h66;
		memory[16'h65a2] <= 8'h62;
		memory[16'h65a3] <= 8'hf5;
		memory[16'h65a4] <= 8'h18;
		memory[16'h65a5] <= 8'h40;
		memory[16'h65a6] <= 8'hb9;
		memory[16'h65a7] <= 8'h76;
		memory[16'h65a8] <= 8'hca;
		memory[16'h65a9] <= 8'hc8;
		memory[16'h65aa] <= 8'h2d;
		memory[16'h65ab] <= 8'h99;
		memory[16'h65ac] <= 8'h91;
		memory[16'h65ad] <= 8'hc9;
		memory[16'h65ae] <= 8'h89;
		memory[16'h65af] <= 8'hff;
		memory[16'h65b0] <= 8'h46;
		memory[16'h65b1] <= 8'hef;
		memory[16'h65b2] <= 8'hd;
		memory[16'h65b3] <= 8'h0;
		memory[16'h65b4] <= 8'h87;
		memory[16'h65b5] <= 8'h4f;
		memory[16'h65b6] <= 8'h6;
		memory[16'h65b7] <= 8'h91;
		memory[16'h65b8] <= 8'he7;
		memory[16'h65b9] <= 8'h8d;
		memory[16'h65ba] <= 8'he3;
		memory[16'h65bb] <= 8'hce;
		memory[16'h65bc] <= 8'ha6;
		memory[16'h65bd] <= 8'hf5;
		memory[16'h65be] <= 8'h4e;
		memory[16'h65bf] <= 8'h54;
		memory[16'h65c0] <= 8'h5c;
		memory[16'h65c1] <= 8'hb1;
		memory[16'h65c2] <= 8'h4a;
		memory[16'h65c3] <= 8'h74;
		memory[16'h65c4] <= 8'hf1;
		memory[16'h65c5] <= 8'h3;
		memory[16'h65c6] <= 8'hea;
		memory[16'h65c7] <= 8'hbb;
		memory[16'h65c8] <= 8'hcb;
		memory[16'h65c9] <= 8'h17;
		memory[16'h65ca] <= 8'h55;
		memory[16'h65cb] <= 8'h5d;
		memory[16'h65cc] <= 8'he0;
		memory[16'h65cd] <= 8'hde;
		memory[16'h65ce] <= 8'h5c;
		memory[16'h65cf] <= 8'h26;
		memory[16'h65d0] <= 8'hcd;
		memory[16'h65d1] <= 8'h6a;
		memory[16'h65d2] <= 8'h26;
		memory[16'h65d3] <= 8'h54;
		memory[16'h65d4] <= 8'hb9;
		memory[16'h65d5] <= 8'h2c;
		memory[16'h65d6] <= 8'he6;
		memory[16'h65d7] <= 8'ha0;
		memory[16'h65d8] <= 8'hb9;
		memory[16'h65d9] <= 8'hc9;
		memory[16'h65da] <= 8'h6f;
		memory[16'h65db] <= 8'h60;
		memory[16'h65dc] <= 8'hbe;
		memory[16'h65dd] <= 8'hbd;
		memory[16'h65de] <= 8'hb4;
		memory[16'h65df] <= 8'h1a;
		memory[16'h65e0] <= 8'h6e;
		memory[16'h65e1] <= 8'hfe;
		memory[16'h65e2] <= 8'h8e;
		memory[16'h65e3] <= 8'h5f;
		memory[16'h65e4] <= 8'h2;
		memory[16'h65e5] <= 8'h78;
		memory[16'h65e6] <= 8'h1b;
		memory[16'h65e7] <= 8'hcd;
		memory[16'h65e8] <= 8'h8f;
		memory[16'h65e9] <= 8'h70;
		memory[16'h65ea] <= 8'h2a;
		memory[16'h65eb] <= 8'h6f;
		memory[16'h65ec] <= 8'h4e;
		memory[16'h65ed] <= 8'h87;
		memory[16'h65ee] <= 8'h96;
		memory[16'h65ef] <= 8'h1b;
		memory[16'h65f0] <= 8'hf1;
		memory[16'h65f1] <= 8'hbc;
		memory[16'h65f2] <= 8'h70;
		memory[16'h65f3] <= 8'haa;
		memory[16'h65f4] <= 8'he9;
		memory[16'h65f5] <= 8'h56;
		memory[16'h65f6] <= 8'h4b;
		memory[16'h65f7] <= 8'ha2;
		memory[16'h65f8] <= 8'h1f;
		memory[16'h65f9] <= 8'hba;
		memory[16'h65fa] <= 8'h2;
		memory[16'h65fb] <= 8'hdd;
		memory[16'h65fc] <= 8'h77;
		memory[16'h65fd] <= 8'hb7;
		memory[16'h65fe] <= 8'hf8;
		memory[16'h65ff] <= 8'he6;
		memory[16'h6600] <= 8'hb5;
		memory[16'h6601] <= 8'h86;
		memory[16'h6602] <= 8'h45;
		memory[16'h6603] <= 8'hb7;
		memory[16'h6604] <= 8'hff;
		memory[16'h6605] <= 8'h60;
		memory[16'h6606] <= 8'h85;
		memory[16'h6607] <= 8'h8e;
		memory[16'h6608] <= 8'hd0;
		memory[16'h6609] <= 8'haf;
		memory[16'h660a] <= 8'hfe;
		memory[16'h660b] <= 8'h1e;
		memory[16'h660c] <= 8'h36;
		memory[16'h660d] <= 8'h94;
		memory[16'h660e] <= 8'h3a;
		memory[16'h660f] <= 8'h27;
		memory[16'h6610] <= 8'h50;
		memory[16'h6611] <= 8'haa;
		memory[16'h6612] <= 8'hd2;
		memory[16'h6613] <= 8'h39;
		memory[16'h6614] <= 8'h0;
		memory[16'h6615] <= 8'h1d;
		memory[16'h6616] <= 8'hdc;
		memory[16'h6617] <= 8'h1f;
		memory[16'h6618] <= 8'hd7;
		memory[16'h6619] <= 8'hde;
		memory[16'h661a] <= 8'hfc;
		memory[16'h661b] <= 8'h4e;
		memory[16'h661c] <= 8'h95;
		memory[16'h661d] <= 8'hf4;
		memory[16'h661e] <= 8'h34;
		memory[16'h661f] <= 8'h4b;
		memory[16'h6620] <= 8'h7b;
		memory[16'h6621] <= 8'h7a;
		memory[16'h6622] <= 8'h2;
		memory[16'h6623] <= 8'h7a;
		memory[16'h6624] <= 8'hda;
		memory[16'h6625] <= 8'h87;
		memory[16'h6626] <= 8'h8;
		memory[16'h6627] <= 8'hab;
		memory[16'h6628] <= 8'h37;
		memory[16'h6629] <= 8'h6;
		memory[16'h662a] <= 8'hc9;
		memory[16'h662b] <= 8'h6d;
		memory[16'h662c] <= 8'h9a;
		memory[16'h662d] <= 8'h3;
		memory[16'h662e] <= 8'h95;
		memory[16'h662f] <= 8'heb;
		memory[16'h6630] <= 8'had;
		memory[16'h6631] <= 8'h67;
		memory[16'h6632] <= 8'h24;
		memory[16'h6633] <= 8'had;
		memory[16'h6634] <= 8'h84;
		memory[16'h6635] <= 8'h0;
		memory[16'h6636] <= 8'hcc;
		memory[16'h6637] <= 8'h5b;
		memory[16'h6638] <= 8'hdf;
		memory[16'h6639] <= 8'hc9;
		memory[16'h663a] <= 8'ha9;
		memory[16'h663b] <= 8'h74;
		memory[16'h663c] <= 8'hbd;
		memory[16'h663d] <= 8'hde;
		memory[16'h663e] <= 8'hbf;
		memory[16'h663f] <= 8'h38;
		memory[16'h6640] <= 8'h58;
		memory[16'h6641] <= 8'hc2;
		memory[16'h6642] <= 8'hb2;
		memory[16'h6643] <= 8'h32;
		memory[16'h6644] <= 8'h49;
		memory[16'h6645] <= 8'hbb;
		memory[16'h6646] <= 8'hdd;
		memory[16'h6647] <= 8'h80;
		memory[16'h6648] <= 8'hc1;
		memory[16'h6649] <= 8'ha7;
		memory[16'h664a] <= 8'hee;
		memory[16'h664b] <= 8'h5c;
		memory[16'h664c] <= 8'haa;
		memory[16'h664d] <= 8'h83;
		memory[16'h664e] <= 8'h47;
		memory[16'h664f] <= 8'h58;
		memory[16'h6650] <= 8'hea;
		memory[16'h6651] <= 8'h6b;
		memory[16'h6652] <= 8'h5;
		memory[16'h6653] <= 8'h6e;
		memory[16'h6654] <= 8'h6c;
		memory[16'h6655] <= 8'hd2;
		memory[16'h6656] <= 8'hc9;
		memory[16'h6657] <= 8'h4b;
		memory[16'h6658] <= 8'h9b;
		memory[16'h6659] <= 8'h72;
		memory[16'h665a] <= 8'hbf;
		memory[16'h665b] <= 8'h58;
		memory[16'h665c] <= 8'h50;
		memory[16'h665d] <= 8'h7f;
		memory[16'h665e] <= 8'h91;
		memory[16'h665f] <= 8'ha8;
		memory[16'h6660] <= 8'h41;
		memory[16'h6661] <= 8'h43;
		memory[16'h6662] <= 8'hdb;
		memory[16'h6663] <= 8'h8a;
		memory[16'h6664] <= 8'hfe;
		memory[16'h6665] <= 8'hb8;
		memory[16'h6666] <= 8'hb;
		memory[16'h6667] <= 8'hc0;
		memory[16'h6668] <= 8'h5f;
		memory[16'h6669] <= 8'hf9;
		memory[16'h666a] <= 8'h1c;
		memory[16'h666b] <= 8'ha;
		memory[16'h666c] <= 8'h7c;
		memory[16'h666d] <= 8'h63;
		memory[16'h666e] <= 8'h62;
		memory[16'h666f] <= 8'h66;
		memory[16'h6670] <= 8'hce;
		memory[16'h6671] <= 8'h67;
		memory[16'h6672] <= 8'hd4;
		memory[16'h6673] <= 8'h3a;
		memory[16'h6674] <= 8'h39;
		memory[16'h6675] <= 8'h9d;
		memory[16'h6676] <= 8'h85;
		memory[16'h6677] <= 8'hd4;
		memory[16'h6678] <= 8'hf;
		memory[16'h6679] <= 8'h45;
		memory[16'h667a] <= 8'h2d;
		memory[16'h667b] <= 8'h60;
		memory[16'h667c] <= 8'hc4;
		memory[16'h667d] <= 8'hbe;
		memory[16'h667e] <= 8'h8;
		memory[16'h667f] <= 8'h5;
		memory[16'h6680] <= 8'h1;
		memory[16'h6681] <= 8'he3;
		memory[16'h6682] <= 8'h8f;
		memory[16'h6683] <= 8'h0;
		memory[16'h6684] <= 8'h9c;
		memory[16'h6685] <= 8'h9a;
		memory[16'h6686] <= 8'hc0;
		memory[16'h6687] <= 8'hfb;
		memory[16'h6688] <= 8'h93;
		memory[16'h6689] <= 8'hdc;
		memory[16'h668a] <= 8'h5;
		memory[16'h668b] <= 8'hf;
		memory[16'h668c] <= 8'h3f;
		memory[16'h668d] <= 8'h67;
		memory[16'h668e] <= 8'h75;
		memory[16'h668f] <= 8'hd;
		memory[16'h6690] <= 8'hcf;
		memory[16'h6691] <= 8'h49;
		memory[16'h6692] <= 8'h48;
		memory[16'h6693] <= 8'h8;
		memory[16'h6694] <= 8'he6;
		memory[16'h6695] <= 8'hcd;
		memory[16'h6696] <= 8'hdd;
		memory[16'h6697] <= 8'hf6;
		memory[16'h6698] <= 8'h12;
		memory[16'h6699] <= 8'ha;
		memory[16'h669a] <= 8'h56;
		memory[16'h669b] <= 8'hd6;
		memory[16'h669c] <= 8'hc8;
		memory[16'h669d] <= 8'h5e;
		memory[16'h669e] <= 8'hdb;
		memory[16'h669f] <= 8'hc9;
		memory[16'h66a0] <= 8'h42;
		memory[16'h66a1] <= 8'h6b;
		memory[16'h66a2] <= 8'hc9;
		memory[16'h66a3] <= 8'hde;
		memory[16'h66a4] <= 8'h5;
		memory[16'h66a5] <= 8'h89;
		memory[16'h66a6] <= 8'hd9;
		memory[16'h66a7] <= 8'h99;
		memory[16'h66a8] <= 8'h65;
		memory[16'h66a9] <= 8'hdf;
		memory[16'h66aa] <= 8'ha8;
		memory[16'h66ab] <= 8'ha4;
		memory[16'h66ac] <= 8'h46;
		memory[16'h66ad] <= 8'h1e;
		memory[16'h66ae] <= 8'hb2;
		memory[16'h66af] <= 8'h15;
		memory[16'h66b0] <= 8'h67;
		memory[16'h66b1] <= 8'hfa;
		memory[16'h66b2] <= 8'h1e;
		memory[16'h66b3] <= 8'h4e;
		memory[16'h66b4] <= 8'hc7;
		memory[16'h66b5] <= 8'hfb;
		memory[16'h66b6] <= 8'h44;
		memory[16'h66b7] <= 8'hda;
		memory[16'h66b8] <= 8'h5;
		memory[16'h66b9] <= 8'h9a;
		memory[16'h66ba] <= 8'hb0;
		memory[16'h66bb] <= 8'hcd;
		memory[16'h66bc] <= 8'hf8;
		memory[16'h66bd] <= 8'h8c;
		memory[16'h66be] <= 8'h96;
		memory[16'h66bf] <= 8'h3a;
		memory[16'h66c0] <= 8'hf7;
		memory[16'h66c1] <= 8'h60;
		memory[16'h66c2] <= 8'h18;
		memory[16'h66c3] <= 8'hfc;
		memory[16'h66c4] <= 8'he9;
		memory[16'h66c5] <= 8'hf2;
		memory[16'h66c6] <= 8'h95;
		memory[16'h66c7] <= 8'h4f;
		memory[16'h66c8] <= 8'hd1;
		memory[16'h66c9] <= 8'h3e;
		memory[16'h66ca] <= 8'hf3;
		memory[16'h66cb] <= 8'h17;
		memory[16'h66cc] <= 8'h5c;
		memory[16'h66cd] <= 8'ha5;
		memory[16'h66ce] <= 8'h2d;
		memory[16'h66cf] <= 8'hc3;
		memory[16'h66d0] <= 8'h9f;
		memory[16'h66d1] <= 8'h4b;
		memory[16'h66d2] <= 8'h11;
		memory[16'h66d3] <= 8'h67;
		memory[16'h66d4] <= 8'h46;
		memory[16'h66d5] <= 8'h55;
		memory[16'h66d6] <= 8'h41;
		memory[16'h66d7] <= 8'h4b;
		memory[16'h66d8] <= 8'hef;
		memory[16'h66d9] <= 8'hf1;
		memory[16'h66da] <= 8'h18;
		memory[16'h66db] <= 8'he8;
		memory[16'h66dc] <= 8'h7d;
		memory[16'h66dd] <= 8'hae;
		memory[16'h66de] <= 8'h22;
		memory[16'h66df] <= 8'h74;
		memory[16'h66e0] <= 8'he;
		memory[16'h66e1] <= 8'h3b;
		memory[16'h66e2] <= 8'h71;
		memory[16'h66e3] <= 8'hf8;
		memory[16'h66e4] <= 8'h2d;
		memory[16'h66e5] <= 8'h6;
		memory[16'h66e6] <= 8'h47;
		memory[16'h66e7] <= 8'hfe;
		memory[16'h66e8] <= 8'h44;
		memory[16'h66e9] <= 8'h3a;
		memory[16'h66ea] <= 8'h15;
		memory[16'h66eb] <= 8'ha0;
		memory[16'h66ec] <= 8'he0;
		memory[16'h66ed] <= 8'h42;
		memory[16'h66ee] <= 8'h64;
		memory[16'h66ef] <= 8'h7f;
		memory[16'h66f0] <= 8'h8d;
		memory[16'h66f1] <= 8'h75;
		memory[16'h66f2] <= 8'he6;
		memory[16'h66f3] <= 8'hd3;
		memory[16'h66f4] <= 8'hcb;
		memory[16'h66f5] <= 8'h27;
		memory[16'h66f6] <= 8'h1e;
		memory[16'h66f7] <= 8'hba;
		memory[16'h66f8] <= 8'h19;
		memory[16'h66f9] <= 8'h36;
		memory[16'h66fa] <= 8'ha2;
		memory[16'h66fb] <= 8'h96;
		memory[16'h66fc] <= 8'he5;
		memory[16'h66fd] <= 8'hc5;
		memory[16'h66fe] <= 8'hb;
		memory[16'h66ff] <= 8'hf3;
		memory[16'h6700] <= 8'h0;
		memory[16'h6701] <= 8'h7c;
		memory[16'h6702] <= 8'heb;
		memory[16'h6703] <= 8'h2d;
		memory[16'h6704] <= 8'h82;
		memory[16'h6705] <= 8'h32;
		memory[16'h6706] <= 8'h2b;
		memory[16'h6707] <= 8'hc7;
		memory[16'h6708] <= 8'h6d;
		memory[16'h6709] <= 8'h40;
		memory[16'h670a] <= 8'h67;
		memory[16'h670b] <= 8'h4d;
		memory[16'h670c] <= 8'h83;
		memory[16'h670d] <= 8'hcb;
		memory[16'h670e] <= 8'hcc;
		memory[16'h670f] <= 8'h10;
		memory[16'h6710] <= 8'h41;
		memory[16'h6711] <= 8'hb3;
		memory[16'h6712] <= 8'he4;
		memory[16'h6713] <= 8'hc;
		memory[16'h6714] <= 8'hda;
		memory[16'h6715] <= 8'h2;
		memory[16'h6716] <= 8'hc6;
		memory[16'h6717] <= 8'hf3;
		memory[16'h6718] <= 8'h39;
		memory[16'h6719] <= 8'h69;
		memory[16'h671a] <= 8'h8a;
		memory[16'h671b] <= 8'h1e;
		memory[16'h671c] <= 8'h2e;
		memory[16'h671d] <= 8'h95;
		memory[16'h671e] <= 8'h11;
		memory[16'h671f] <= 8'h2e;
		memory[16'h6720] <= 8'h11;
		memory[16'h6721] <= 8'hfd;
		memory[16'h6722] <= 8'h5b;
		memory[16'h6723] <= 8'h93;
		memory[16'h6724] <= 8'h2f;
		memory[16'h6725] <= 8'h86;
		memory[16'h6726] <= 8'h5a;
		memory[16'h6727] <= 8'h9c;
		memory[16'h6728] <= 8'hc6;
		memory[16'h6729] <= 8'hc2;
		memory[16'h672a] <= 8'he9;
		memory[16'h672b] <= 8'h49;
		memory[16'h672c] <= 8'h8d;
		memory[16'h672d] <= 8'hb6;
		memory[16'h672e] <= 8'h5a;
		memory[16'h672f] <= 8'hce;
		memory[16'h6730] <= 8'h69;
		memory[16'h6731] <= 8'h3e;
		memory[16'h6732] <= 8'hda;
		memory[16'h6733] <= 8'h43;
		memory[16'h6734] <= 8'h40;
		memory[16'h6735] <= 8'ha1;
		memory[16'h6736] <= 8'h37;
		memory[16'h6737] <= 8'h79;
		memory[16'h6738] <= 8'ha;
		memory[16'h6739] <= 8'hc1;
		memory[16'h673a] <= 8'h97;
		memory[16'h673b] <= 8'h38;
		memory[16'h673c] <= 8'h56;
		memory[16'h673d] <= 8'ha9;
		memory[16'h673e] <= 8'h66;
		memory[16'h673f] <= 8'h67;
		memory[16'h6740] <= 8'ha6;
		memory[16'h6741] <= 8'hc1;
		memory[16'h6742] <= 8'hfa;
		memory[16'h6743] <= 8'hd5;
		memory[16'h6744] <= 8'h47;
		memory[16'h6745] <= 8'h55;
		memory[16'h6746] <= 8'h72;
		memory[16'h6747] <= 8'hd;
		memory[16'h6748] <= 8'h17;
		memory[16'h6749] <= 8'h5b;
		memory[16'h674a] <= 8'h57;
		memory[16'h674b] <= 8'ha4;
		memory[16'h674c] <= 8'h11;
		memory[16'h674d] <= 8'hb1;
		memory[16'h674e] <= 8'h73;
		memory[16'h674f] <= 8'h7a;
		memory[16'h6750] <= 8'hef;
		memory[16'h6751] <= 8'h4d;
		memory[16'h6752] <= 8'hbe;
		memory[16'h6753] <= 8'h2f;
		memory[16'h6754] <= 8'hee;
		memory[16'h6755] <= 8'hf5;
		memory[16'h6756] <= 8'ha9;
		memory[16'h6757] <= 8'hf8;
		memory[16'h6758] <= 8'hb6;
		memory[16'h6759] <= 8'h40;
		memory[16'h675a] <= 8'h30;
		memory[16'h675b] <= 8'hc;
		memory[16'h675c] <= 8'he9;
		memory[16'h675d] <= 8'h96;
		memory[16'h675e] <= 8'h73;
		memory[16'h675f] <= 8'h8f;
		memory[16'h6760] <= 8'h57;
		memory[16'h6761] <= 8'h6d;
		memory[16'h6762] <= 8'h65;
		memory[16'h6763] <= 8'h9e;
		memory[16'h6764] <= 8'hc2;
		memory[16'h6765] <= 8'hd7;
		memory[16'h6766] <= 8'hac;
		memory[16'h6767] <= 8'hd9;
		memory[16'h6768] <= 8'h32;
		memory[16'h6769] <= 8'h3;
		memory[16'h676a] <= 8'h7e;
		memory[16'h676b] <= 8'h44;
		memory[16'h676c] <= 8'hb4;
		memory[16'h676d] <= 8'hf1;
		memory[16'h676e] <= 8'hbe;
		memory[16'h676f] <= 8'ha3;
		memory[16'h6770] <= 8'h3e;
		memory[16'h6771] <= 8'h7c;
		memory[16'h6772] <= 8'hd2;
		memory[16'h6773] <= 8'h2d;
		memory[16'h6774] <= 8'h71;
		memory[16'h6775] <= 8'h7b;
		memory[16'h6776] <= 8'h25;
		memory[16'h6777] <= 8'h27;
		memory[16'h6778] <= 8'hbc;
		memory[16'h6779] <= 8'h56;
		memory[16'h677a] <= 8'h33;
		memory[16'h677b] <= 8'ha5;
		memory[16'h677c] <= 8'hec;
		memory[16'h677d] <= 8'ha6;
		memory[16'h677e] <= 8'h35;
		memory[16'h677f] <= 8'h44;
		memory[16'h6780] <= 8'h14;
		memory[16'h6781] <= 8'h9a;
		memory[16'h6782] <= 8'he2;
		memory[16'h6783] <= 8'hd6;
		memory[16'h6784] <= 8'h71;
		memory[16'h6785] <= 8'h8e;
		memory[16'h6786] <= 8'hb0;
		memory[16'h6787] <= 8'ha3;
		memory[16'h6788] <= 8'h91;
		memory[16'h6789] <= 8'h2e;
		memory[16'h678a] <= 8'he7;
		memory[16'h678b] <= 8'h45;
		memory[16'h678c] <= 8'h1f;
		memory[16'h678d] <= 8'ha6;
		memory[16'h678e] <= 8'he8;
		memory[16'h678f] <= 8'h5d;
		memory[16'h6790] <= 8'h22;
		memory[16'h6791] <= 8'hbb;
		memory[16'h6792] <= 8'h8a;
		memory[16'h6793] <= 8'h94;
		memory[16'h6794] <= 8'h36;
		memory[16'h6795] <= 8'hb0;
		memory[16'h6796] <= 8'hbb;
		memory[16'h6797] <= 8'hf2;
		memory[16'h6798] <= 8'h6;
		memory[16'h6799] <= 8'hef;
		memory[16'h679a] <= 8'h98;
		memory[16'h679b] <= 8'hf2;
		memory[16'h679c] <= 8'h95;
		memory[16'h679d] <= 8'hcd;
		memory[16'h679e] <= 8'h36;
		memory[16'h679f] <= 8'ha9;
		memory[16'h67a0] <= 8'h67;
		memory[16'h67a1] <= 8'h19;
		memory[16'h67a2] <= 8'h80;
		memory[16'h67a3] <= 8'hd8;
		memory[16'h67a4] <= 8'ha7;
		memory[16'h67a5] <= 8'h30;
		memory[16'h67a6] <= 8'h7b;
		memory[16'h67a7] <= 8'h39;
		memory[16'h67a8] <= 8'h5e;
		memory[16'h67a9] <= 8'h63;
		memory[16'h67aa] <= 8'h7e;
		memory[16'h67ab] <= 8'h7d;
		memory[16'h67ac] <= 8'h9;
		memory[16'h67ad] <= 8'h67;
		memory[16'h67ae] <= 8'hda;
		memory[16'h67af] <= 8'h2b;
		memory[16'h67b0] <= 8'h22;
		memory[16'h67b1] <= 8'h65;
		memory[16'h67b2] <= 8'hbf;
		memory[16'h67b3] <= 8'h58;
		memory[16'h67b4] <= 8'h15;
		memory[16'h67b5] <= 8'h7b;
		memory[16'h67b6] <= 8'h4b;
		memory[16'h67b7] <= 8'h1b;
		memory[16'h67b8] <= 8'h6a;
		memory[16'h67b9] <= 8'he3;
		memory[16'h67ba] <= 8'hd;
		memory[16'h67bb] <= 8'hff;
		memory[16'h67bc] <= 8'hb0;
		memory[16'h67bd] <= 8'h44;
		memory[16'h67be] <= 8'ha9;
		memory[16'h67bf] <= 8'h17;
		memory[16'h67c0] <= 8'h5d;
		memory[16'h67c1] <= 8'h29;
		memory[16'h67c2] <= 8'hef;
		memory[16'h67c3] <= 8'h4;
		memory[16'h67c4] <= 8'h59;
		memory[16'h67c5] <= 8'h6a;
		memory[16'h67c6] <= 8'h3d;
		memory[16'h67c7] <= 8'hb7;
		memory[16'h67c8] <= 8'hcd;
		memory[16'h67c9] <= 8'hbc;
		memory[16'h67ca] <= 8'h34;
		memory[16'h67cb] <= 8'hd6;
		memory[16'h67cc] <= 8'h23;
		memory[16'h67cd] <= 8'he;
		memory[16'h67ce] <= 8'h2;
		memory[16'h67cf] <= 8'h45;
		memory[16'h67d0] <= 8'h73;
		memory[16'h67d1] <= 8'hc1;
		memory[16'h67d2] <= 8'h9d;
		memory[16'h67d3] <= 8'h88;
		memory[16'h67d4] <= 8'h3c;
		memory[16'h67d5] <= 8'he8;
		memory[16'h67d6] <= 8'ha3;
		memory[16'h67d7] <= 8'ha6;
		memory[16'h67d8] <= 8'hcb;
		memory[16'h67d9] <= 8'hb1;
		memory[16'h67da] <= 8'ha6;
		memory[16'h67db] <= 8'h7b;
		memory[16'h67dc] <= 8'hf5;
		memory[16'h67dd] <= 8'h4f;
		memory[16'h67de] <= 8'h92;
		memory[16'h67df] <= 8'h52;
		memory[16'h67e0] <= 8'h78;
		memory[16'h67e1] <= 8'h81;
		memory[16'h67e2] <= 8'h56;
		memory[16'h67e3] <= 8'hd1;
		memory[16'h67e4] <= 8'hec;
		memory[16'h67e5] <= 8'h94;
		memory[16'h67e6] <= 8'h88;
		memory[16'h67e7] <= 8'hb9;
		memory[16'h67e8] <= 8'h50;
		memory[16'h67e9] <= 8'hbc;
		memory[16'h67ea] <= 8'h90;
		memory[16'h67eb] <= 8'h73;
		memory[16'h67ec] <= 8'hca;
		memory[16'h67ed] <= 8'h92;
		memory[16'h67ee] <= 8'hb8;
		memory[16'h67ef] <= 8'h3e;
		memory[16'h67f0] <= 8'h53;
		memory[16'h67f1] <= 8'h55;
		memory[16'h67f2] <= 8'hc6;
		memory[16'h67f3] <= 8'h90;
		memory[16'h67f4] <= 8'h3e;
		memory[16'h67f5] <= 8'h6a;
		memory[16'h67f6] <= 8'h36;
		memory[16'h67f7] <= 8'h9;
		memory[16'h67f8] <= 8'h1b;
		memory[16'h67f9] <= 8'hdc;
		memory[16'h67fa] <= 8'h85;
		memory[16'h67fb] <= 8'h10;
		memory[16'h67fc] <= 8'h2b;
		memory[16'h67fd] <= 8'h17;
		memory[16'h67fe] <= 8'h62;
		memory[16'h67ff] <= 8'ha3;
		memory[16'h6800] <= 8'h99;
		memory[16'h6801] <= 8'hb8;
		memory[16'h6802] <= 8'h74;
		memory[16'h6803] <= 8'h85;
		memory[16'h6804] <= 8'h4c;
		memory[16'h6805] <= 8'hfc;
		memory[16'h6806] <= 8'h3e;
		memory[16'h6807] <= 8'h9c;
		memory[16'h6808] <= 8'hb8;
		memory[16'h6809] <= 8'hce;
		memory[16'h680a] <= 8'hf;
		memory[16'h680b] <= 8'h83;
		memory[16'h680c] <= 8'h60;
		memory[16'h680d] <= 8'hc7;
		memory[16'h680e] <= 8'hc1;
		memory[16'h680f] <= 8'hb4;
		memory[16'h6810] <= 8'h1d;
		memory[16'h6811] <= 8'h87;
		memory[16'h6812] <= 8'h44;
		memory[16'h6813] <= 8'h5b;
		memory[16'h6814] <= 8'hf1;
		memory[16'h6815] <= 8'h7a;
		memory[16'h6816] <= 8'h64;
		memory[16'h6817] <= 8'hc;
		memory[16'h6818] <= 8'h57;
		memory[16'h6819] <= 8'he9;
		memory[16'h681a] <= 8'h1c;
		memory[16'h681b] <= 8'h82;
		memory[16'h681c] <= 8'h1;
		memory[16'h681d] <= 8'h7e;
		memory[16'h681e] <= 8'h26;
		memory[16'h681f] <= 8'h9a;
		memory[16'h6820] <= 8'h37;
		memory[16'h6821] <= 8'h9a;
		memory[16'h6822] <= 8'h1f;
		memory[16'h6823] <= 8'h83;
		memory[16'h6824] <= 8'h97;
		memory[16'h6825] <= 8'h5d;
		memory[16'h6826] <= 8'h20;
		memory[16'h6827] <= 8'h4f;
		memory[16'h6828] <= 8'h2c;
		memory[16'h6829] <= 8'h2f;
		memory[16'h682a] <= 8'hd2;
		memory[16'h682b] <= 8'h8c;
		memory[16'h682c] <= 8'hf7;
		memory[16'h682d] <= 8'h93;
		memory[16'h682e] <= 8'h40;
		memory[16'h682f] <= 8'h14;
		memory[16'h6830] <= 8'h1b;
		memory[16'h6831] <= 8'h84;
		memory[16'h6832] <= 8'h6f;
		memory[16'h6833] <= 8'hc;
		memory[16'h6834] <= 8'hff;
		memory[16'h6835] <= 8'hd3;
		memory[16'h6836] <= 8'h19;
		memory[16'h6837] <= 8'h56;
		memory[16'h6838] <= 8'hbd;
		memory[16'h6839] <= 8'h35;
		memory[16'h683a] <= 8'hd8;
		memory[16'h683b] <= 8'hbe;
		memory[16'h683c] <= 8'hb4;
		memory[16'h683d] <= 8'hfe;
		memory[16'h683e] <= 8'h58;
		memory[16'h683f] <= 8'heb;
		memory[16'h6840] <= 8'h99;
		memory[16'h6841] <= 8'h77;
		memory[16'h6842] <= 8'h6e;
		memory[16'h6843] <= 8'h30;
		memory[16'h6844] <= 8'hd4;
		memory[16'h6845] <= 8'h8e;
		memory[16'h6846] <= 8'h7f;
		memory[16'h6847] <= 8'h0;
		memory[16'h6848] <= 8'hbe;
		memory[16'h6849] <= 8'h52;
		memory[16'h684a] <= 8'h8d;
		memory[16'h684b] <= 8'hb5;
		memory[16'h684c] <= 8'he5;
		memory[16'h684d] <= 8'hcd;
		memory[16'h684e] <= 8'hc9;
		memory[16'h684f] <= 8'h0;
		memory[16'h6850] <= 8'h52;
		memory[16'h6851] <= 8'h38;
		memory[16'h6852] <= 8'hd;
		memory[16'h6853] <= 8'h51;
		memory[16'h6854] <= 8'hb;
		memory[16'h6855] <= 8'h26;
		memory[16'h6856] <= 8'ha7;
		memory[16'h6857] <= 8'hc8;
		memory[16'h6858] <= 8'h5b;
		memory[16'h6859] <= 8'h7f;
		memory[16'h685a] <= 8'h86;
		memory[16'h685b] <= 8'hf;
		memory[16'h685c] <= 8'h7e;
		memory[16'h685d] <= 8'hde;
		memory[16'h685e] <= 8'hfa;
		memory[16'h685f] <= 8'h17;
		memory[16'h6860] <= 8'h55;
		memory[16'h6861] <= 8'h69;
		memory[16'h6862] <= 8'h47;
		memory[16'h6863] <= 8'h2a;
		memory[16'h6864] <= 8'hf7;
		memory[16'h6865] <= 8'hc6;
		memory[16'h6866] <= 8'h2a;
		memory[16'h6867] <= 8'hb5;
		memory[16'h6868] <= 8'h18;
		memory[16'h6869] <= 8'hb7;
		memory[16'h686a] <= 8'h6a;
		memory[16'h686b] <= 8'hfe;
		memory[16'h686c] <= 8'h85;
		memory[16'h686d] <= 8'h33;
		memory[16'h686e] <= 8'hfe;
		memory[16'h686f] <= 8'hd7;
		memory[16'h6870] <= 8'h6b;
		memory[16'h6871] <= 8'hb;
		memory[16'h6872] <= 8'h28;
		memory[16'h6873] <= 8'h77;
		memory[16'h6874] <= 8'h31;
		memory[16'h6875] <= 8'hcf;
		memory[16'h6876] <= 8'h3f;
		memory[16'h6877] <= 8'h8d;
		memory[16'h6878] <= 8'h4e;
		memory[16'h6879] <= 8'hc6;
		memory[16'h687a] <= 8'h9c;
		memory[16'h687b] <= 8'hcc;
		memory[16'h687c] <= 8'ha4;
		memory[16'h687d] <= 8'h97;
		memory[16'h687e] <= 8'he3;
		memory[16'h687f] <= 8'hfa;
		memory[16'h6880] <= 8'h0;
		memory[16'h6881] <= 8'h2a;
		memory[16'h6882] <= 8'h24;
		memory[16'h6883] <= 8'hf7;
		memory[16'h6884] <= 8'hf1;
		memory[16'h6885] <= 8'h4e;
		memory[16'h6886] <= 8'had;
		memory[16'h6887] <= 8'h9;
		memory[16'h6888] <= 8'h6;
		memory[16'h6889] <= 8'h17;
		memory[16'h688a] <= 8'h7;
		memory[16'h688b] <= 8'h8b;
		memory[16'h688c] <= 8'h4b;
		memory[16'h688d] <= 8'h6;
		memory[16'h688e] <= 8'h62;
		memory[16'h688f] <= 8'hb6;
		memory[16'h6890] <= 8'h11;
		memory[16'h6891] <= 8'h8a;
		memory[16'h6892] <= 8'h2d;
		memory[16'h6893] <= 8'h43;
		memory[16'h6894] <= 8'h59;
		memory[16'h6895] <= 8'h6d;
		memory[16'h6896] <= 8'hd0;
		memory[16'h6897] <= 8'ha7;
		memory[16'h6898] <= 8'h33;
		memory[16'h6899] <= 8'h6c;
		memory[16'h689a] <= 8'h74;
		memory[16'h689b] <= 8'hd7;
		memory[16'h689c] <= 8'h3;
		memory[16'h689d] <= 8'h57;
		memory[16'h689e] <= 8'hd1;
		memory[16'h689f] <= 8'h3;
		memory[16'h68a0] <= 8'h82;
		memory[16'h68a1] <= 8'hf5;
		memory[16'h68a2] <= 8'hfb;
		memory[16'h68a3] <= 8'h73;
		memory[16'h68a4] <= 8'h44;
		memory[16'h68a5] <= 8'ha8;
		memory[16'h68a6] <= 8'h7c;
		memory[16'h68a7] <= 8'h4a;
		memory[16'h68a8] <= 8'hbf;
		memory[16'h68a9] <= 8'h84;
		memory[16'h68aa] <= 8'hd5;
		memory[16'h68ab] <= 8'ha;
		memory[16'h68ac] <= 8'h8a;
		memory[16'h68ad] <= 8'h37;
		memory[16'h68ae] <= 8'hc1;
		memory[16'h68af] <= 8'h9b;
		memory[16'h68b0] <= 8'hc1;
		memory[16'h68b1] <= 8'hee;
		memory[16'h68b2] <= 8'hde;
		memory[16'h68b3] <= 8'h1a;
		memory[16'h68b4] <= 8'h5b;
		memory[16'h68b5] <= 8'hae;
		memory[16'h68b6] <= 8'hc1;
		memory[16'h68b7] <= 8'h8e;
		memory[16'h68b8] <= 8'h1b;
		memory[16'h68b9] <= 8'h35;
		memory[16'h68ba] <= 8'h66;
		memory[16'h68bb] <= 8'h1e;
		memory[16'h68bc] <= 8'h8d;
		memory[16'h68bd] <= 8'h37;
		memory[16'h68be] <= 8'h22;
		memory[16'h68bf] <= 8'hf;
		memory[16'h68c0] <= 8'h2d;
		memory[16'h68c1] <= 8'h1d;
		memory[16'h68c2] <= 8'h82;
		memory[16'h68c3] <= 8'h71;
		memory[16'h68c4] <= 8'hc5;
		memory[16'h68c5] <= 8'hfe;
		memory[16'h68c6] <= 8'hbb;
		memory[16'h68c7] <= 8'h84;
		memory[16'h68c8] <= 8'h82;
		memory[16'h68c9] <= 8'h90;
		memory[16'h68ca] <= 8'h8f;
		memory[16'h68cb] <= 8'hc;
		memory[16'h68cc] <= 8'hc7;
		memory[16'h68cd] <= 8'h50;
		memory[16'h68ce] <= 8'ha8;
		memory[16'h68cf] <= 8'h88;
		memory[16'h68d0] <= 8'h3e;
		memory[16'h68d1] <= 8'h86;
		memory[16'h68d2] <= 8'ha2;
		memory[16'h68d3] <= 8'h9a;
		memory[16'h68d4] <= 8'h35;
		memory[16'h68d5] <= 8'h63;
		memory[16'h68d6] <= 8'h28;
		memory[16'h68d7] <= 8'h50;
		memory[16'h68d8] <= 8'h99;
		memory[16'h68d9] <= 8'h8e;
		memory[16'h68da] <= 8'h6e;
		memory[16'h68db] <= 8'h26;
		memory[16'h68dc] <= 8'hc6;
		memory[16'h68dd] <= 8'h90;
		memory[16'h68de] <= 8'h35;
		memory[16'h68df] <= 8'hf3;
		memory[16'h68e0] <= 8'had;
		memory[16'h68e1] <= 8'hb7;
		memory[16'h68e2] <= 8'h64;
		memory[16'h68e3] <= 8'h72;
		memory[16'h68e4] <= 8'hb5;
		memory[16'h68e5] <= 8'h1f;
		memory[16'h68e6] <= 8'hf7;
		memory[16'h68e7] <= 8'h38;
		memory[16'h68e8] <= 8'haf;
		memory[16'h68e9] <= 8'h86;
		memory[16'h68ea] <= 8'h44;
		memory[16'h68eb] <= 8'h76;
		memory[16'h68ec] <= 8'hd6;
		memory[16'h68ed] <= 8'hec;
		memory[16'h68ee] <= 8'hfe;
		memory[16'h68ef] <= 8'h14;
		memory[16'h68f0] <= 8'h73;
		memory[16'h68f1] <= 8'ha0;
		memory[16'h68f2] <= 8'hae;
		memory[16'h68f3] <= 8'ha8;
		memory[16'h68f4] <= 8'h3;
		memory[16'h68f5] <= 8'hd7;
		memory[16'h68f6] <= 8'hf8;
		memory[16'h68f7] <= 8'h9c;
		memory[16'h68f8] <= 8'h65;
		memory[16'h68f9] <= 8'h66;
		memory[16'h68fa] <= 8'hc2;
		memory[16'h68fb] <= 8'h2b;
		memory[16'h68fc] <= 8'hf7;
		memory[16'h68fd] <= 8'hf7;
		memory[16'h68fe] <= 8'h1e;
		memory[16'h68ff] <= 8'ha4;
		memory[16'h6900] <= 8'hae;
		memory[16'h6901] <= 8'h82;
		memory[16'h6902] <= 8'h17;
		memory[16'h6903] <= 8'h64;
		memory[16'h6904] <= 8'ha1;
		memory[16'h6905] <= 8'he;
		memory[16'h6906] <= 8'h9c;
		memory[16'h6907] <= 8'h50;
		memory[16'h6908] <= 8'h94;
		memory[16'h6909] <= 8'he0;
		memory[16'h690a] <= 8'hc6;
		memory[16'h690b] <= 8'h6a;
		memory[16'h690c] <= 8'hcd;
		memory[16'h690d] <= 8'hc4;
		memory[16'h690e] <= 8'h7e;
		memory[16'h690f] <= 8'h40;
		memory[16'h6910] <= 8'h64;
		memory[16'h6911] <= 8'h2d;
		memory[16'h6912] <= 8'he8;
		memory[16'h6913] <= 8'h68;
		memory[16'h6914] <= 8'h4;
		memory[16'h6915] <= 8'he0;
		memory[16'h6916] <= 8'h4;
		memory[16'h6917] <= 8'h69;
		memory[16'h6918] <= 8'h46;
		memory[16'h6919] <= 8'hc7;
		memory[16'h691a] <= 8'h95;
		memory[16'h691b] <= 8'h3d;
		memory[16'h691c] <= 8'hbe;
		memory[16'h691d] <= 8'hb3;
		memory[16'h691e] <= 8'he2;
		memory[16'h691f] <= 8'h6d;
		memory[16'h6920] <= 8'h36;
		memory[16'h6921] <= 8'hf9;
		memory[16'h6922] <= 8'hd1;
		memory[16'h6923] <= 8'hd7;
		memory[16'h6924] <= 8'h7;
		memory[16'h6925] <= 8'h6d;
		memory[16'h6926] <= 8'h28;
		memory[16'h6927] <= 8'h9b;
		memory[16'h6928] <= 8'h4d;
		memory[16'h6929] <= 8'hee;
		memory[16'h692a] <= 8'h5;
		memory[16'h692b] <= 8'h1a;
		memory[16'h692c] <= 8'hb3;
		memory[16'h692d] <= 8'h83;
		memory[16'h692e] <= 8'h5a;
		memory[16'h692f] <= 8'h17;
		memory[16'h6930] <= 8'hb0;
		memory[16'h6931] <= 8'h42;
		memory[16'h6932] <= 8'h7f;
		memory[16'h6933] <= 8'hb4;
		memory[16'h6934] <= 8'h22;
		memory[16'h6935] <= 8'h84;
		memory[16'h6936] <= 8'h1e;
		memory[16'h6937] <= 8'h69;
		memory[16'h6938] <= 8'h4b;
		memory[16'h6939] <= 8'hb3;
		memory[16'h693a] <= 8'ha6;
		memory[16'h693b] <= 8'h9;
		memory[16'h693c] <= 8'h66;
		memory[16'h693d] <= 8'h88;
		memory[16'h693e] <= 8'h76;
		memory[16'h693f] <= 8'h9c;
		memory[16'h6940] <= 8'h81;
		memory[16'h6941] <= 8'h47;
		memory[16'h6942] <= 8'h74;
		memory[16'h6943] <= 8'h88;
		memory[16'h6944] <= 8'hb4;
		memory[16'h6945] <= 8'h9c;
		memory[16'h6946] <= 8'h23;
		memory[16'h6947] <= 8'h2;
		memory[16'h6948] <= 8'h8a;
		memory[16'h6949] <= 8'h28;
		memory[16'h694a] <= 8'h1c;
		memory[16'h694b] <= 8'h3d;
		memory[16'h694c] <= 8'hac;
		memory[16'h694d] <= 8'h77;
		memory[16'h694e] <= 8'h55;
		memory[16'h694f] <= 8'h5c;
		memory[16'h6950] <= 8'hb9;
		memory[16'h6951] <= 8'hd4;
		memory[16'h6952] <= 8'h11;
		memory[16'h6953] <= 8'hdc;
		memory[16'h6954] <= 8'h58;
		memory[16'h6955] <= 8'h2f;
		memory[16'h6956] <= 8'h45;
		memory[16'h6957] <= 8'ha3;
		memory[16'h6958] <= 8'he2;
		memory[16'h6959] <= 8'heb;
		memory[16'h695a] <= 8'had;
		memory[16'h695b] <= 8'h48;
		memory[16'h695c] <= 8'h74;
		memory[16'h695d] <= 8'h23;
		memory[16'h695e] <= 8'he5;
		memory[16'h695f] <= 8'hf5;
		memory[16'h6960] <= 8'h6b;
		memory[16'h6961] <= 8'h59;
		memory[16'h6962] <= 8'h7e;
		memory[16'h6963] <= 8'h1f;
		memory[16'h6964] <= 8'hf5;
		memory[16'h6965] <= 8'ha1;
		memory[16'h6966] <= 8'h21;
		memory[16'h6967] <= 8'h7f;
		memory[16'h6968] <= 8'hca;
		memory[16'h6969] <= 8'h3e;
		memory[16'h696a] <= 8'hbd;
		memory[16'h696b] <= 8'h76;
		memory[16'h696c] <= 8'hb5;
		memory[16'h696d] <= 8'h12;
		memory[16'h696e] <= 8'hd2;
		memory[16'h696f] <= 8'h6e;
		memory[16'h6970] <= 8'he6;
		memory[16'h6971] <= 8'he3;
		memory[16'h6972] <= 8'h4a;
		memory[16'h6973] <= 8'h3f;
		memory[16'h6974] <= 8'h12;
		memory[16'h6975] <= 8'h8f;
		memory[16'h6976] <= 8'he2;
		memory[16'h6977] <= 8'hf4;
		memory[16'h6978] <= 8'h7b;
		memory[16'h6979] <= 8'h8f;
		memory[16'h697a] <= 8'h3d;
		memory[16'h697b] <= 8'hef;
		memory[16'h697c] <= 8'hb3;
		memory[16'h697d] <= 8'h22;
		memory[16'h697e] <= 8'he4;
		memory[16'h697f] <= 8'h1e;
		memory[16'h6980] <= 8'h7b;
		memory[16'h6981] <= 8'h62;
		memory[16'h6982] <= 8'h3d;
		memory[16'h6983] <= 8'h70;
		memory[16'h6984] <= 8'h4;
		memory[16'h6985] <= 8'h5f;
		memory[16'h6986] <= 8'hef;
		memory[16'h6987] <= 8'hce;
		memory[16'h6988] <= 8'h9d;
		memory[16'h6989] <= 8'hac;
		memory[16'h698a] <= 8'h44;
		memory[16'h698b] <= 8'h52;
		memory[16'h698c] <= 8'hbe;
		memory[16'h698d] <= 8'h16;
		memory[16'h698e] <= 8'hc0;
		memory[16'h698f] <= 8'ha5;
		memory[16'h6990] <= 8'hfa;
		memory[16'h6991] <= 8'hb;
		memory[16'h6992] <= 8'he4;
		memory[16'h6993] <= 8'hc;
		memory[16'h6994] <= 8'h9a;
		memory[16'h6995] <= 8'hc6;
		memory[16'h6996] <= 8'h1;
		memory[16'h6997] <= 8'h15;
		memory[16'h6998] <= 8'h56;
		memory[16'h6999] <= 8'h3e;
		memory[16'h699a] <= 8'h4;
		memory[16'h699b] <= 8'h9;
		memory[16'h699c] <= 8'h60;
		memory[16'h699d] <= 8'he9;
		memory[16'h699e] <= 8'h27;
		memory[16'h699f] <= 8'hdb;
		memory[16'h69a0] <= 8'h4b;
		memory[16'h69a1] <= 8'h64;
		memory[16'h69a2] <= 8'h4b;
		memory[16'h69a3] <= 8'h4f;
		memory[16'h69a4] <= 8'hc3;
		memory[16'h69a5] <= 8'h3a;
		memory[16'h69a6] <= 8'h1d;
		memory[16'h69a7] <= 8'h60;
		memory[16'h69a8] <= 8'he7;
		memory[16'h69a9] <= 8'h61;
		memory[16'h69aa] <= 8'hb2;
		memory[16'h69ab] <= 8'ha5;
		memory[16'h69ac] <= 8'h78;
		memory[16'h69ad] <= 8'h73;
		memory[16'h69ae] <= 8'h4a;
		memory[16'h69af] <= 8'h72;
		memory[16'h69b0] <= 8'h7e;
		memory[16'h69b1] <= 8'h2e;
		memory[16'h69b2] <= 8'h7e;
		memory[16'h69b3] <= 8'h18;
		memory[16'h69b4] <= 8'hf5;
		memory[16'h69b5] <= 8'h7f;
		memory[16'h69b6] <= 8'h2e;
		memory[16'h69b7] <= 8'h4b;
		memory[16'h69b8] <= 8'hbd;
		memory[16'h69b9] <= 8'h32;
		memory[16'h69ba] <= 8'h54;
		memory[16'h69bb] <= 8'h1d;
		memory[16'h69bc] <= 8'h1b;
		memory[16'h69bd] <= 8'h7b;
		memory[16'h69be] <= 8'hf8;
		memory[16'h69bf] <= 8'h67;
		memory[16'h69c0] <= 8'hdf;
		memory[16'h69c1] <= 8'h43;
		memory[16'h69c2] <= 8'hb6;
		memory[16'h69c3] <= 8'ha3;
		memory[16'h69c4] <= 8'h7e;
		memory[16'h69c5] <= 8'hd4;
		memory[16'h69c6] <= 8'h3;
		memory[16'h69c7] <= 8'h65;
		memory[16'h69c8] <= 8'h35;
		memory[16'h69c9] <= 8'hb6;
		memory[16'h69ca] <= 8'ha;
		memory[16'h69cb] <= 8'had;
		memory[16'h69cc] <= 8'h29;
		memory[16'h69cd] <= 8'h55;
		memory[16'h69ce] <= 8'h1f;
		memory[16'h69cf] <= 8'ha7;
		memory[16'h69d0] <= 8'h83;
		memory[16'h69d1] <= 8'h9e;
		memory[16'h69d2] <= 8'hbf;
		memory[16'h69d3] <= 8'h78;
		memory[16'h69d4] <= 8'h1d;
		memory[16'h69d5] <= 8'hed;
		memory[16'h69d6] <= 8'hc3;
		memory[16'h69d7] <= 8'hdb;
		memory[16'h69d8] <= 8'h20;
		memory[16'h69d9] <= 8'h17;
		memory[16'h69da] <= 8'hf8;
		memory[16'h69db] <= 8'h3b;
		memory[16'h69dc] <= 8'h92;
		memory[16'h69dd] <= 8'hf1;
		memory[16'h69de] <= 8'ha2;
		memory[16'h69df] <= 8'h72;
		memory[16'h69e0] <= 8'h34;
		memory[16'h69e1] <= 8'h59;
		memory[16'h69e2] <= 8'h15;
		memory[16'h69e3] <= 8'hb2;
		memory[16'h69e4] <= 8'h2d;
		memory[16'h69e5] <= 8'h18;
		memory[16'h69e6] <= 8'h17;
		memory[16'h69e7] <= 8'h62;
		memory[16'h69e8] <= 8'hce;
		memory[16'h69e9] <= 8'h22;
		memory[16'h69ea] <= 8'h10;
		memory[16'h69eb] <= 8'hf7;
		memory[16'h69ec] <= 8'h77;
		memory[16'h69ed] <= 8'h2f;
		memory[16'h69ee] <= 8'h9e;
		memory[16'h69ef] <= 8'hfa;
		memory[16'h69f0] <= 8'hcd;
		memory[16'h69f1] <= 8'h5e;
		memory[16'h69f2] <= 8'h73;
		memory[16'h69f3] <= 8'heb;
		memory[16'h69f4] <= 8'h4b;
		memory[16'h69f5] <= 8'h36;
		memory[16'h69f6] <= 8'hc6;
		memory[16'h69f7] <= 8'h6b;
		memory[16'h69f8] <= 8'h4e;
		memory[16'h69f9] <= 8'hbe;
		memory[16'h69fa] <= 8'ha7;
		memory[16'h69fb] <= 8'he0;
		memory[16'h69fc] <= 8'haf;
		memory[16'h69fd] <= 8'h49;
		memory[16'h69fe] <= 8'h52;
		memory[16'h69ff] <= 8'he4;
		memory[16'h6a00] <= 8'ha2;
		memory[16'h6a01] <= 8'h67;
		memory[16'h6a02] <= 8'h96;
		memory[16'h6a03] <= 8'hcf;
		memory[16'h6a04] <= 8'h80;
		memory[16'h6a05] <= 8'hae;
		memory[16'h6a06] <= 8'h32;
		memory[16'h6a07] <= 8'h4e;
		memory[16'h6a08] <= 8'hd0;
		memory[16'h6a09] <= 8'h42;
		memory[16'h6a0a] <= 8'h46;
		memory[16'h6a0b] <= 8'h47;
		memory[16'h6a0c] <= 8'h71;
		memory[16'h6a0d] <= 8'he4;
		memory[16'h6a0e] <= 8'h41;
		memory[16'h6a0f] <= 8'h3f;
		memory[16'h6a10] <= 8'h42;
		memory[16'h6a11] <= 8'hb4;
		memory[16'h6a12] <= 8'h2a;
		memory[16'h6a13] <= 8'h8e;
		memory[16'h6a14] <= 8'heb;
		memory[16'h6a15] <= 8'hf0;
		memory[16'h6a16] <= 8'hf9;
		memory[16'h6a17] <= 8'h39;
		memory[16'h6a18] <= 8'hae;
		memory[16'h6a19] <= 8'ha0;
		memory[16'h6a1a] <= 8'h19;
		memory[16'h6a1b] <= 8'h5e;
		memory[16'h6a1c] <= 8'hea;
		memory[16'h6a1d] <= 8'h6c;
		memory[16'h6a1e] <= 8'h42;
		memory[16'h6a1f] <= 8'h8c;
		memory[16'h6a20] <= 8'hd3;
		memory[16'h6a21] <= 8'hd8;
		memory[16'h6a22] <= 8'h5c;
		memory[16'h6a23] <= 8'h53;
		memory[16'h6a24] <= 8'h86;
		memory[16'h6a25] <= 8'h8e;
		memory[16'h6a26] <= 8'ha2;
		memory[16'h6a27] <= 8'h56;
		memory[16'h6a28] <= 8'hd0;
		memory[16'h6a29] <= 8'he8;
		memory[16'h6a2a] <= 8'h9d;
		memory[16'h6a2b] <= 8'h41;
		memory[16'h6a2c] <= 8'hcc;
		memory[16'h6a2d] <= 8'hdf;
		memory[16'h6a2e] <= 8'h80;
		memory[16'h6a2f] <= 8'hf;
		memory[16'h6a30] <= 8'h93;
		memory[16'h6a31] <= 8'haa;
		memory[16'h6a32] <= 8'h9d;
		memory[16'h6a33] <= 8'h7e;
		memory[16'h6a34] <= 8'h9a;
		memory[16'h6a35] <= 8'h96;
		memory[16'h6a36] <= 8'hb7;
		memory[16'h6a37] <= 8'h49;
		memory[16'h6a38] <= 8'h37;
		memory[16'h6a39] <= 8'hd1;
		memory[16'h6a3a] <= 8'ha7;
		memory[16'h6a3b] <= 8'h21;
		memory[16'h6a3c] <= 8'h3d;
		memory[16'h6a3d] <= 8'he9;
		memory[16'h6a3e] <= 8'had;
		memory[16'h6a3f] <= 8'h10;
		memory[16'h6a40] <= 8'hc1;
		memory[16'h6a41] <= 8'h9;
		memory[16'h6a42] <= 8'h64;
		memory[16'h6a43] <= 8'h48;
		memory[16'h6a44] <= 8'h97;
		memory[16'h6a45] <= 8'h6;
		memory[16'h6a46] <= 8'h9e;
		memory[16'h6a47] <= 8'h67;
		memory[16'h6a48] <= 8'hee;
		memory[16'h6a49] <= 8'h3c;
		memory[16'h6a4a] <= 8'ha9;
		memory[16'h6a4b] <= 8'hba;
		memory[16'h6a4c] <= 8'h1b;
		memory[16'h6a4d] <= 8'h29;
		memory[16'h6a4e] <= 8'hc9;
		memory[16'h6a4f] <= 8'hae;
		memory[16'h6a50] <= 8'hd4;
		memory[16'h6a51] <= 8'h66;
		memory[16'h6a52] <= 8'h2d;
		memory[16'h6a53] <= 8'h6e;
		memory[16'h6a54] <= 8'hfd;
		memory[16'h6a55] <= 8'he4;
		memory[16'h6a56] <= 8'hb7;
		memory[16'h6a57] <= 8'h34;
		memory[16'h6a58] <= 8'hb5;
		memory[16'h6a59] <= 8'h5e;
		memory[16'h6a5a] <= 8'h55;
		memory[16'h6a5b] <= 8'hf2;
		memory[16'h6a5c] <= 8'h47;
		memory[16'h6a5d] <= 8'h2;
		memory[16'h6a5e] <= 8'h3;
		memory[16'h6a5f] <= 8'h9;
		memory[16'h6a60] <= 8'hc;
		memory[16'h6a61] <= 8'h67;
		memory[16'h6a62] <= 8'h51;
		memory[16'h6a63] <= 8'ha3;
		memory[16'h6a64] <= 8'h6d;
		memory[16'h6a65] <= 8'hef;
		memory[16'h6a66] <= 8'hb;
		memory[16'h6a67] <= 8'h5b;
		memory[16'h6a68] <= 8'h2b;
		memory[16'h6a69] <= 8'hb4;
		memory[16'h6a6a] <= 8'h15;
		memory[16'h6a6b] <= 8'h46;
		memory[16'h6a6c] <= 8'hdd;
		memory[16'h6a6d] <= 8'hdf;
		memory[16'h6a6e] <= 8'hf5;
		memory[16'h6a6f] <= 8'hb1;
		memory[16'h6a70] <= 8'h45;
		memory[16'h6a71] <= 8'h22;
		memory[16'h6a72] <= 8'h20;
		memory[16'h6a73] <= 8'h42;
		memory[16'h6a74] <= 8'h6;
		memory[16'h6a75] <= 8'hd7;
		memory[16'h6a76] <= 8'h76;
		memory[16'h6a77] <= 8'hbc;
		memory[16'h6a78] <= 8'h36;
		memory[16'h6a79] <= 8'hcb;
		memory[16'h6a7a] <= 8'hae;
		memory[16'h6a7b] <= 8'h7d;
		memory[16'h6a7c] <= 8'hce;
		memory[16'h6a7d] <= 8'hb1;
		memory[16'h6a7e] <= 8'h86;
		memory[16'h6a7f] <= 8'hda;
		memory[16'h6a80] <= 8'h18;
		memory[16'h6a81] <= 8'hd7;
		memory[16'h6a82] <= 8'h7d;
		memory[16'h6a83] <= 8'h85;
		memory[16'h6a84] <= 8'hc7;
		memory[16'h6a85] <= 8'h88;
		memory[16'h6a86] <= 8'he0;
		memory[16'h6a87] <= 8'hf2;
		memory[16'h6a88] <= 8'h3c;
		memory[16'h6a89] <= 8'hf6;
		memory[16'h6a8a] <= 8'h39;
		memory[16'h6a8b] <= 8'h1a;
		memory[16'h6a8c] <= 8'hd5;
		memory[16'h6a8d] <= 8'h2e;
		memory[16'h6a8e] <= 8'hcb;
		memory[16'h6a8f] <= 8'h1a;
		memory[16'h6a90] <= 8'h50;
		memory[16'h6a91] <= 8'heb;
		memory[16'h6a92] <= 8'h5d;
		memory[16'h6a93] <= 8'h56;
		memory[16'h6a94] <= 8'hc3;
		memory[16'h6a95] <= 8'hd3;
		memory[16'h6a96] <= 8'h12;
		memory[16'h6a97] <= 8'hf9;
		memory[16'h6a98] <= 8'h9f;
		memory[16'h6a99] <= 8'hc1;
		memory[16'h6a9a] <= 8'h76;
		memory[16'h6a9b] <= 8'h6d;
		memory[16'h6a9c] <= 8'h72;
		memory[16'h6a9d] <= 8'hfd;
		memory[16'h6a9e] <= 8'h47;
		memory[16'h6a9f] <= 8'h8b;
		memory[16'h6aa0] <= 8'hd4;
		memory[16'h6aa1] <= 8'hc4;
		memory[16'h6aa2] <= 8'h10;
		memory[16'h6aa3] <= 8'h9b;
		memory[16'h6aa4] <= 8'h4d;
		memory[16'h6aa5] <= 8'hf1;
		memory[16'h6aa6] <= 8'h8e;
		memory[16'h6aa7] <= 8'h89;
		memory[16'h6aa8] <= 8'he7;
		memory[16'h6aa9] <= 8'hc7;
		memory[16'h6aaa] <= 8'ha3;
		memory[16'h6aab] <= 8'hbc;
		memory[16'h6aac] <= 8'hf5;
		memory[16'h6aad] <= 8'h6f;
		memory[16'h6aae] <= 8'hd6;
		memory[16'h6aaf] <= 8'h45;
		memory[16'h6ab0] <= 8'h5a;
		memory[16'h6ab1] <= 8'h33;
		memory[16'h6ab2] <= 8'h9b;
		memory[16'h6ab3] <= 8'h1d;
		memory[16'h6ab4] <= 8'h7;
		memory[16'h6ab5] <= 8'hae;
		memory[16'h6ab6] <= 8'h16;
		memory[16'h6ab7] <= 8'ha6;
		memory[16'h6ab8] <= 8'h6f;
		memory[16'h6ab9] <= 8'h8d;
		memory[16'h6aba] <= 8'h13;
		memory[16'h6abb] <= 8'he1;
		memory[16'h6abc] <= 8'h8a;
		memory[16'h6abd] <= 8'h5a;
		memory[16'h6abe] <= 8'h6c;
		memory[16'h6abf] <= 8'h5e;
		memory[16'h6ac0] <= 8'h1e;
		memory[16'h6ac1] <= 8'h7d;
		memory[16'h6ac2] <= 8'hfa;
		memory[16'h6ac3] <= 8'h6b;
		memory[16'h6ac4] <= 8'h6e;
		memory[16'h6ac5] <= 8'h88;
		memory[16'h6ac6] <= 8'hf5;
		memory[16'h6ac7] <= 8'h55;
		memory[16'h6ac8] <= 8'h4f;
		memory[16'h6ac9] <= 8'h98;
		memory[16'h6aca] <= 8'h11;
		memory[16'h6acb] <= 8'h44;
		memory[16'h6acc] <= 8'h7;
		memory[16'h6acd] <= 8'he7;
		memory[16'h6ace] <= 8'h89;
		memory[16'h6acf] <= 8'h62;
		memory[16'h6ad0] <= 8'h1b;
		memory[16'h6ad1] <= 8'h24;
		memory[16'h6ad2] <= 8'h7f;
		memory[16'h6ad3] <= 8'h22;
		memory[16'h6ad4] <= 8'hd2;
		memory[16'h6ad5] <= 8'h96;
		memory[16'h6ad6] <= 8'hc8;
		memory[16'h6ad7] <= 8'h41;
		memory[16'h6ad8] <= 8'h23;
		memory[16'h6ad9] <= 8'hdb;
		memory[16'h6ada] <= 8'h23;
		memory[16'h6adb] <= 8'had;
		memory[16'h6adc] <= 8'h35;
		memory[16'h6add] <= 8'h8f;
		memory[16'h6ade] <= 8'hb;
		memory[16'h6adf] <= 8'h53;
		memory[16'h6ae0] <= 8'hc;
		memory[16'h6ae1] <= 8'h5;
		memory[16'h6ae2] <= 8'hbf;
		memory[16'h6ae3] <= 8'h7a;
		memory[16'h6ae4] <= 8'h8d;
		memory[16'h6ae5] <= 8'hb4;
		memory[16'h6ae6] <= 8'hcf;
		memory[16'h6ae7] <= 8'hdc;
		memory[16'h6ae8] <= 8'h4c;
		memory[16'h6ae9] <= 8'he0;
		memory[16'h6aea] <= 8'h20;
		memory[16'h6aeb] <= 8'h54;
		memory[16'h6aec] <= 8'hc8;
		memory[16'h6aed] <= 8'ha9;
		memory[16'h6aee] <= 8'hb6;
		memory[16'h6aef] <= 8'he3;
		memory[16'h6af0] <= 8'hce;
		memory[16'h6af1] <= 8'h35;
		memory[16'h6af2] <= 8'h5;
		memory[16'h6af3] <= 8'ha0;
		memory[16'h6af4] <= 8'hcb;
		memory[16'h6af5] <= 8'hcd;
		memory[16'h6af6] <= 8'he2;
		memory[16'h6af7] <= 8'hee;
		memory[16'h6af8] <= 8'ha8;
		memory[16'h6af9] <= 8'h5;
		memory[16'h6afa] <= 8'h9b;
		memory[16'h6afb] <= 8'hdd;
		memory[16'h6afc] <= 8'h94;
		memory[16'h6afd] <= 8'ha7;
		memory[16'h6afe] <= 8'h30;
		memory[16'h6aff] <= 8'ha1;
		memory[16'h6b00] <= 8'hac;
		memory[16'h6b01] <= 8'hef;
		memory[16'h6b02] <= 8'h1b;
		memory[16'h6b03] <= 8'h3a;
		memory[16'h6b04] <= 8'ha3;
		memory[16'h6b05] <= 8'heb;
		memory[16'h6b06] <= 8'h16;
		memory[16'h6b07] <= 8'hf0;
		memory[16'h6b08] <= 8'hcb;
		memory[16'h6b09] <= 8'h37;
		memory[16'h6b0a] <= 8'h44;
		memory[16'h6b0b] <= 8'h93;
		memory[16'h6b0c] <= 8'he0;
		memory[16'h6b0d] <= 8'hfa;
		memory[16'h6b0e] <= 8'h76;
		memory[16'h6b0f] <= 8'hae;
		memory[16'h6b10] <= 8'h2f;
		memory[16'h6b11] <= 8'h7b;
		memory[16'h6b12] <= 8'h4f;
		memory[16'h6b13] <= 8'hfb;
		memory[16'h6b14] <= 8'h48;
		memory[16'h6b15] <= 8'h31;
		memory[16'h6b16] <= 8'he9;
		memory[16'h6b17] <= 8'hf0;
		memory[16'h6b18] <= 8'h36;
		memory[16'h6b19] <= 8'h85;
		memory[16'h6b1a] <= 8'hcd;
		memory[16'h6b1b] <= 8'hca;
		memory[16'h6b1c] <= 8'h2c;
		memory[16'h6b1d] <= 8'hfe;
		memory[16'h6b1e] <= 8'h6b;
		memory[16'h6b1f] <= 8'hd8;
		memory[16'h6b20] <= 8'hed;
		memory[16'h6b21] <= 8'h87;
		memory[16'h6b22] <= 8'h12;
		memory[16'h6b23] <= 8'h91;
		memory[16'h6b24] <= 8'h72;
		memory[16'h6b25] <= 8'h29;
		memory[16'h6b26] <= 8'h81;
		memory[16'h6b27] <= 8'h3d;
		memory[16'h6b28] <= 8'h60;
		memory[16'h6b29] <= 8'hc5;
		memory[16'h6b2a] <= 8'hd1;
		memory[16'h6b2b] <= 8'h40;
		memory[16'h6b2c] <= 8'hbf;
		memory[16'h6b2d] <= 8'h47;
		memory[16'h6b2e] <= 8'hef;
		memory[16'h6b2f] <= 8'hee;
		memory[16'h6b30] <= 8'hc3;
		memory[16'h6b31] <= 8'h3e;
		memory[16'h6b32] <= 8'he9;
		memory[16'h6b33] <= 8'hb;
		memory[16'h6b34] <= 8'h6f;
		memory[16'h6b35] <= 8'hd3;
		memory[16'h6b36] <= 8'hfc;
		memory[16'h6b37] <= 8'ha5;
		memory[16'h6b38] <= 8'h58;
		memory[16'h6b39] <= 8'hc9;
		memory[16'h6b3a] <= 8'h6f;
		memory[16'h6b3b] <= 8'h84;
		memory[16'h6b3c] <= 8'hc7;
		memory[16'h6b3d] <= 8'hdb;
		memory[16'h6b3e] <= 8'h5c;
		memory[16'h6b3f] <= 8'hb5;
		memory[16'h6b40] <= 8'h62;
		memory[16'h6b41] <= 8'h6f;
		memory[16'h6b42] <= 8'h46;
		memory[16'h6b43] <= 8'hd4;
		memory[16'h6b44] <= 8'h98;
		memory[16'h6b45] <= 8'hc7;
		memory[16'h6b46] <= 8'h11;
		memory[16'h6b47] <= 8'hf8;
		memory[16'h6b48] <= 8'h8c;
		memory[16'h6b49] <= 8'he2;
		memory[16'h6b4a] <= 8'h38;
		memory[16'h6b4b] <= 8'h4b;
		memory[16'h6b4c] <= 8'h2a;
		memory[16'h6b4d] <= 8'h27;
		memory[16'h6b4e] <= 8'h39;
		memory[16'h6b4f] <= 8'hed;
		memory[16'h6b50] <= 8'h65;
		memory[16'h6b51] <= 8'h23;
		memory[16'h6b52] <= 8'hf8;
		memory[16'h6b53] <= 8'hd4;
		memory[16'h6b54] <= 8'hf6;
		memory[16'h6b55] <= 8'hf4;
		memory[16'h6b56] <= 8'h79;
		memory[16'h6b57] <= 8'h4e;
		memory[16'h6b58] <= 8'hbe;
		memory[16'h6b59] <= 8'he9;
		memory[16'h6b5a] <= 8'hd2;
		memory[16'h6b5b] <= 8'h85;
		memory[16'h6b5c] <= 8'hc4;
		memory[16'h6b5d] <= 8'h2e;
		memory[16'h6b5e] <= 8'h3a;
		memory[16'h6b5f] <= 8'h26;
		memory[16'h6b60] <= 8'h9d;
		memory[16'h6b61] <= 8'h80;
		memory[16'h6b62] <= 8'hfa;
		memory[16'h6b63] <= 8'h35;
		memory[16'h6b64] <= 8'h47;
		memory[16'h6b65] <= 8'hb;
		memory[16'h6b66] <= 8'h2d;
		memory[16'h6b67] <= 8'hd3;
		memory[16'h6b68] <= 8'hee;
		memory[16'h6b69] <= 8'h66;
		memory[16'h6b6a] <= 8'h1e;
		memory[16'h6b6b] <= 8'h18;
		memory[16'h6b6c] <= 8'h8d;
		memory[16'h6b6d] <= 8'h58;
		memory[16'h6b6e] <= 8'h5;
		memory[16'h6b6f] <= 8'hf3;
		memory[16'h6b70] <= 8'h7b;
		memory[16'h6b71] <= 8'hfd;
		memory[16'h6b72] <= 8'hc7;
		memory[16'h6b73] <= 8'h71;
		memory[16'h6b74] <= 8'hf2;
		memory[16'h6b75] <= 8'h41;
		memory[16'h6b76] <= 8'hbf;
		memory[16'h6b77] <= 8'hb0;
		memory[16'h6b78] <= 8'h2a;
		memory[16'h6b79] <= 8'h91;
		memory[16'h6b7a] <= 8'h35;
		memory[16'h6b7b] <= 8'hee;
		memory[16'h6b7c] <= 8'hbf;
		memory[16'h6b7d] <= 8'h70;
		memory[16'h6b7e] <= 8'h14;
		memory[16'h6b7f] <= 8'h5d;
		memory[16'h6b80] <= 8'hf0;
		memory[16'h6b81] <= 8'he;
		memory[16'h6b82] <= 8'h92;
		memory[16'h6b83] <= 8'h38;
		memory[16'h6b84] <= 8'h19;
		memory[16'h6b85] <= 8'hc0;
		memory[16'h6b86] <= 8'hb;
		memory[16'h6b87] <= 8'h7;
		memory[16'h6b88] <= 8'h26;
		memory[16'h6b89] <= 8'h2a;
		memory[16'h6b8a] <= 8'h1f;
		memory[16'h6b8b] <= 8'hb3;
		memory[16'h6b8c] <= 8'h82;
		memory[16'h6b8d] <= 8'h24;
		memory[16'h6b8e] <= 8'ha6;
		memory[16'h6b8f] <= 8'hfd;
		memory[16'h6b90] <= 8'h22;
		memory[16'h6b91] <= 8'h6e;
		memory[16'h6b92] <= 8'h6e;
		memory[16'h6b93] <= 8'h14;
		memory[16'h6b94] <= 8'haf;
		memory[16'h6b95] <= 8'h2d;
		memory[16'h6b96] <= 8'hc4;
		memory[16'h6b97] <= 8'hd9;
		memory[16'h6b98] <= 8'hbe;
		memory[16'h6b99] <= 8'hf9;
		memory[16'h6b9a] <= 8'hc7;
		memory[16'h6b9b] <= 8'h7d;
		memory[16'h6b9c] <= 8'h69;
		memory[16'h6b9d] <= 8'hdb;
		memory[16'h6b9e] <= 8'hda;
		memory[16'h6b9f] <= 8'h5a;
		memory[16'h6ba0] <= 8'he9;
		memory[16'h6ba1] <= 8'h6d;
		memory[16'h6ba2] <= 8'h92;
		memory[16'h6ba3] <= 8'h2;
		memory[16'h6ba4] <= 8'h2d;
		memory[16'h6ba5] <= 8'h9d;
		memory[16'h6ba6] <= 8'ha;
		memory[16'h6ba7] <= 8'h53;
		memory[16'h6ba8] <= 8'hc7;
		memory[16'h6ba9] <= 8'h29;
		memory[16'h6baa] <= 8'h6;
		memory[16'h6bab] <= 8'h49;
		memory[16'h6bac] <= 8'h4e;
		memory[16'h6bad] <= 8'had;
		memory[16'h6bae] <= 8'h46;
		memory[16'h6baf] <= 8'h70;
		memory[16'h6bb0] <= 8'h1b;
		memory[16'h6bb1] <= 8'hb4;
		memory[16'h6bb2] <= 8'h84;
		memory[16'h6bb3] <= 8'hca;
		memory[16'h6bb4] <= 8'he1;
		memory[16'h6bb5] <= 8'h48;
		memory[16'h6bb6] <= 8'ha3;
		memory[16'h6bb7] <= 8'h9f;
		memory[16'h6bb8] <= 8'h41;
		memory[16'h6bb9] <= 8'h6a;
		memory[16'h6bba] <= 8'h1d;
		memory[16'h6bbb] <= 8'hab;
		memory[16'h6bbc] <= 8'h45;
		memory[16'h6bbd] <= 8'hf7;
		memory[16'h6bbe] <= 8'h5;
		memory[16'h6bbf] <= 8'h2e;
		memory[16'h6bc0] <= 8'h64;
		memory[16'h6bc1] <= 8'h97;
		memory[16'h6bc2] <= 8'h30;
		memory[16'h6bc3] <= 8'h91;
		memory[16'h6bc4] <= 8'h34;
		memory[16'h6bc5] <= 8'h3a;
		memory[16'h6bc6] <= 8'he4;
		memory[16'h6bc7] <= 8'hfc;
		memory[16'h6bc8] <= 8'h64;
		memory[16'h6bc9] <= 8'heb;
		memory[16'h6bca] <= 8'h45;
		memory[16'h6bcb] <= 8'hb2;
		memory[16'h6bcc] <= 8'h98;
		memory[16'h6bcd] <= 8'h8c;
		memory[16'h6bce] <= 8'h22;
		memory[16'h6bcf] <= 8'hb3;
		memory[16'h6bd0] <= 8'h40;
		memory[16'h6bd1] <= 8'ha6;
		memory[16'h6bd2] <= 8'h7d;
		memory[16'h6bd3] <= 8'h22;
		memory[16'h6bd4] <= 8'hee;
		memory[16'h6bd5] <= 8'h20;
		memory[16'h6bd6] <= 8'hc1;
		memory[16'h6bd7] <= 8'h2f;
		memory[16'h6bd8] <= 8'h8a;
		memory[16'h6bd9] <= 8'hde;
		memory[16'h6bda] <= 8'hda;
		memory[16'h6bdb] <= 8'hcf;
		memory[16'h6bdc] <= 8'hd6;
		memory[16'h6bdd] <= 8'hdf;
		memory[16'h6bde] <= 8'hfd;
		memory[16'h6bdf] <= 8'h3a;
		memory[16'h6be0] <= 8'h76;
		memory[16'h6be1] <= 8'h2d;
		memory[16'h6be2] <= 8'hcc;
		memory[16'h6be3] <= 8'hab;
		memory[16'h6be4] <= 8'h68;
		memory[16'h6be5] <= 8'hb0;
		memory[16'h6be6] <= 8'ha7;
		memory[16'h6be7] <= 8'hcc;
		memory[16'h6be8] <= 8'h9b;
		memory[16'h6be9] <= 8'hec;
		memory[16'h6bea] <= 8'h7e;
		memory[16'h6beb] <= 8'h33;
		memory[16'h6bec] <= 8'h78;
		memory[16'h6bed] <= 8'ha0;
		memory[16'h6bee] <= 8'he6;
		memory[16'h6bef] <= 8'hb9;
		memory[16'h6bf0] <= 8'h46;
		memory[16'h6bf1] <= 8'h63;
		memory[16'h6bf2] <= 8'hdb;
		memory[16'h6bf3] <= 8'h34;
		memory[16'h6bf4] <= 8'h83;
		memory[16'h6bf5] <= 8'h9c;
		memory[16'h6bf6] <= 8'h63;
		memory[16'h6bf7] <= 8'hd;
		memory[16'h6bf8] <= 8'h7b;
		memory[16'h6bf9] <= 8'h3e;
		memory[16'h6bfa] <= 8'hdc;
		memory[16'h6bfb] <= 8'h51;
		memory[16'h6bfc] <= 8'h1d;
		memory[16'h6bfd] <= 8'hd9;
		memory[16'h6bfe] <= 8'h8b;
		memory[16'h6bff] <= 8'h94;
		memory[16'h6c00] <= 8'h7;
		memory[16'h6c01] <= 8'h57;
		memory[16'h6c02] <= 8'h3f;
		memory[16'h6c03] <= 8'h6f;
		memory[16'h6c04] <= 8'h8;
		memory[16'h6c05] <= 8'he6;
		memory[16'h6c06] <= 8'h3b;
		memory[16'h6c07] <= 8'ha3;
		memory[16'h6c08] <= 8'hd2;
		memory[16'h6c09] <= 8'hb9;
		memory[16'h6c0a] <= 8'hd7;
		memory[16'h6c0b] <= 8'h4b;
		memory[16'h6c0c] <= 8'h59;
		memory[16'h6c0d] <= 8'hbd;
		memory[16'h6c0e] <= 8'h4;
		memory[16'h6c0f] <= 8'h9f;
		memory[16'h6c10] <= 8'h21;
		memory[16'h6c11] <= 8'hdf;
		memory[16'h6c12] <= 8'hd3;
		memory[16'h6c13] <= 8'ha4;
		memory[16'h6c14] <= 8'h7b;
		memory[16'h6c15] <= 8'h36;
		memory[16'h6c16] <= 8'hb2;
		memory[16'h6c17] <= 8'hf6;
		memory[16'h6c18] <= 8'h74;
		memory[16'h6c19] <= 8'h8e;
		memory[16'h6c1a] <= 8'h47;
		memory[16'h6c1b] <= 8'h92;
		memory[16'h6c1c] <= 8'h68;
		memory[16'h6c1d] <= 8'hd3;
		memory[16'h6c1e] <= 8'h26;
		memory[16'h6c1f] <= 8'h6f;
		memory[16'h6c20] <= 8'h2a;
		memory[16'h6c21] <= 8'h65;
		memory[16'h6c22] <= 8'hde;
		memory[16'h6c23] <= 8'h32;
		memory[16'h6c24] <= 8'h4b;
		memory[16'h6c25] <= 8'h19;
		memory[16'h6c26] <= 8'hd6;
		memory[16'h6c27] <= 8'h1d;
		memory[16'h6c28] <= 8'hd2;
		memory[16'h6c29] <= 8'had;
		memory[16'h6c2a] <= 8'h68;
		memory[16'h6c2b] <= 8'h2b;
		memory[16'h6c2c] <= 8'h6a;
		memory[16'h6c2d] <= 8'h6c;
		memory[16'h6c2e] <= 8'hca;
		memory[16'h6c2f] <= 8'h8b;
		memory[16'h6c30] <= 8'h4b;
		memory[16'h6c31] <= 8'h9d;
		memory[16'h6c32] <= 8'h30;
		memory[16'h6c33] <= 8'hc7;
		memory[16'h6c34] <= 8'hd3;
		memory[16'h6c35] <= 8'he2;
		memory[16'h6c36] <= 8'hbd;
		memory[16'h6c37] <= 8'h48;
		memory[16'h6c38] <= 8'h70;
		memory[16'h6c39] <= 8'h5;
		memory[16'h6c3a] <= 8'hda;
		memory[16'h6c3b] <= 8'hd8;
		memory[16'h6c3c] <= 8'hd8;
		memory[16'h6c3d] <= 8'h0;
		memory[16'h6c3e] <= 8'h47;
		memory[16'h6c3f] <= 8'h2;
		memory[16'h6c40] <= 8'h65;
		memory[16'h6c41] <= 8'h25;
		memory[16'h6c42] <= 8'h35;
		memory[16'h6c43] <= 8'hb0;
		memory[16'h6c44] <= 8'h3e;
		memory[16'h6c45] <= 8'hb;
		memory[16'h6c46] <= 8'hcd;
		memory[16'h6c47] <= 8'h10;
		memory[16'h6c48] <= 8'hb8;
		memory[16'h6c49] <= 8'h36;
		memory[16'h6c4a] <= 8'h3b;
		memory[16'h6c4b] <= 8'h22;
		memory[16'h6c4c] <= 8'ha2;
		memory[16'h6c4d] <= 8'h5;
		memory[16'h6c4e] <= 8'hae;
		memory[16'h6c4f] <= 8'hee;
		memory[16'h6c50] <= 8'ha2;
		memory[16'h6c51] <= 8'hde;
		memory[16'h6c52] <= 8'hb5;
		memory[16'h6c53] <= 8'h76;
		memory[16'h6c54] <= 8'hc0;
		memory[16'h6c55] <= 8'h72;
		memory[16'h6c56] <= 8'hbe;
		memory[16'h6c57] <= 8'h30;
		memory[16'h6c58] <= 8'h77;
		memory[16'h6c59] <= 8'h98;
		memory[16'h6c5a] <= 8'h9;
		memory[16'h6c5b] <= 8'h4f;
		memory[16'h6c5c] <= 8'h98;
		memory[16'h6c5d] <= 8'h50;
		memory[16'h6c5e] <= 8'h52;
		memory[16'h6c5f] <= 8'hfd;
		memory[16'h6c60] <= 8'h76;
		memory[16'h6c61] <= 8'h87;
		memory[16'h6c62] <= 8'had;
		memory[16'h6c63] <= 8'hb4;
		memory[16'h6c64] <= 8'h92;
		memory[16'h6c65] <= 8'h7a;
		memory[16'h6c66] <= 8'hc5;
		memory[16'h6c67] <= 8'h4a;
		memory[16'h6c68] <= 8'hb0;
		memory[16'h6c69] <= 8'h0;
		memory[16'h6c6a] <= 8'h6c;
		memory[16'h6c6b] <= 8'h53;
		memory[16'h6c6c] <= 8'h6;
		memory[16'h6c6d] <= 8'h1a;
		memory[16'h6c6e] <= 8'h41;
		memory[16'h6c6f] <= 8'ha8;
		memory[16'h6c70] <= 8'hf8;
		memory[16'h6c71] <= 8'hf6;
		memory[16'h6c72] <= 8'h1e;
		memory[16'h6c73] <= 8'hb8;
		memory[16'h6c74] <= 8'h68;
		memory[16'h6c75] <= 8'hdc;
		memory[16'h6c76] <= 8'he9;
		memory[16'h6c77] <= 8'he0;
		memory[16'h6c78] <= 8'h74;
		memory[16'h6c79] <= 8'hf2;
		memory[16'h6c7a] <= 8'h2f;
		memory[16'h6c7b] <= 8'hc;
		memory[16'h6c7c] <= 8'h42;
		memory[16'h6c7d] <= 8'h81;
		memory[16'h6c7e] <= 8'h9;
		memory[16'h6c7f] <= 8'hb8;
		memory[16'h6c80] <= 8'h8;
		memory[16'h6c81] <= 8'hb6;
		memory[16'h6c82] <= 8'h6d;
		memory[16'h6c83] <= 8'h9a;
		memory[16'h6c84] <= 8'h31;
		memory[16'h6c85] <= 8'h32;
		memory[16'h6c86] <= 8'he4;
		memory[16'h6c87] <= 8'he1;
		memory[16'h6c88] <= 8'h32;
		memory[16'h6c89] <= 8'h51;
		memory[16'h6c8a] <= 8'h34;
		memory[16'h6c8b] <= 8'h38;
		memory[16'h6c8c] <= 8'h6b;
		memory[16'h6c8d] <= 8'h75;
		memory[16'h6c8e] <= 8'he1;
		memory[16'h6c8f] <= 8'h64;
		memory[16'h6c90] <= 8'h6b;
		memory[16'h6c91] <= 8'hff;
		memory[16'h6c92] <= 8'h1c;
		memory[16'h6c93] <= 8'hd4;
		memory[16'h6c94] <= 8'hdc;
		memory[16'h6c95] <= 8'h5;
		memory[16'h6c96] <= 8'hb4;
		memory[16'h6c97] <= 8'h50;
		memory[16'h6c98] <= 8'hf7;
		memory[16'h6c99] <= 8'he3;
		memory[16'h6c9a] <= 8'h5d;
		memory[16'h6c9b] <= 8'h3a;
		memory[16'h6c9c] <= 8'h65;
		memory[16'h6c9d] <= 8'h66;
		memory[16'h6c9e] <= 8'hf2;
		memory[16'h6c9f] <= 8'h6d;
		memory[16'h6ca0] <= 8'h1d;
		memory[16'h6ca1] <= 8'h5f;
		memory[16'h6ca2] <= 8'h8;
		memory[16'h6ca3] <= 8'h4e;
		memory[16'h6ca4] <= 8'h91;
		memory[16'h6ca5] <= 8'hec;
		memory[16'h6ca6] <= 8'h2f;
		memory[16'h6ca7] <= 8'hc4;
		memory[16'h6ca8] <= 8'h3d;
		memory[16'h6ca9] <= 8'h64;
		memory[16'h6caa] <= 8'hfc;
		memory[16'h6cab] <= 8'ha9;
		memory[16'h6cac] <= 8'hd9;
		memory[16'h6cad] <= 8'hdd;
		memory[16'h6cae] <= 8'hd;
		memory[16'h6caf] <= 8'h45;
		memory[16'h6cb0] <= 8'hdd;
		memory[16'h6cb1] <= 8'h29;
		memory[16'h6cb2] <= 8'h19;
		memory[16'h6cb3] <= 8'hb9;
		memory[16'h6cb4] <= 8'h2f;
		memory[16'h6cb5] <= 8'hcd;
		memory[16'h6cb6] <= 8'h9;
		memory[16'h6cb7] <= 8'h26;
		memory[16'h6cb8] <= 8'hb0;
		memory[16'h6cb9] <= 8'h66;
		memory[16'h6cba] <= 8'h60;
		memory[16'h6cbb] <= 8'h15;
		memory[16'h6cbc] <= 8'hcd;
		memory[16'h6cbd] <= 8'h53;
		memory[16'h6cbe] <= 8'h83;
		memory[16'h6cbf] <= 8'hea;
		memory[16'h6cc0] <= 8'hb2;
		memory[16'h6cc1] <= 8'h8b;
		memory[16'h6cc2] <= 8'h38;
		memory[16'h6cc3] <= 8'h44;
		memory[16'h6cc4] <= 8'h77;
		memory[16'h6cc5] <= 8'h67;
		memory[16'h6cc6] <= 8'h8;
		memory[16'h6cc7] <= 8'hb5;
		memory[16'h6cc8] <= 8'hcb;
		memory[16'h6cc9] <= 8'h4;
		memory[16'h6cca] <= 8'h5e;
		memory[16'h6ccb] <= 8'ha5;
		memory[16'h6ccc] <= 8'he2;
		memory[16'h6ccd] <= 8'h6b;
		memory[16'h6cce] <= 8'hea;
		memory[16'h6ccf] <= 8'hbf;
		memory[16'h6cd0] <= 8'h94;
		memory[16'h6cd1] <= 8'h3;
		memory[16'h6cd2] <= 8'h78;
		memory[16'h6cd3] <= 8'hc3;
		memory[16'h6cd4] <= 8'hd0;
		memory[16'h6cd5] <= 8'h81;
		memory[16'h6cd6] <= 8'hea;
		memory[16'h6cd7] <= 8'h80;
		memory[16'h6cd8] <= 8'he8;
		memory[16'h6cd9] <= 8'h4a;
		memory[16'h6cda] <= 8'h96;
		memory[16'h6cdb] <= 8'hb5;
		memory[16'h6cdc] <= 8'h9d;
		memory[16'h6cdd] <= 8'h19;
		memory[16'h6cde] <= 8'h9f;
		memory[16'h6cdf] <= 8'h50;
		memory[16'h6ce0] <= 8'ha4;
		memory[16'h6ce1] <= 8'hd7;
		memory[16'h6ce2] <= 8'h94;
		memory[16'h6ce3] <= 8'h1b;
		memory[16'h6ce4] <= 8'h3e;
		memory[16'h6ce5] <= 8'h9c;
		memory[16'h6ce6] <= 8'hd0;
		memory[16'h6ce7] <= 8'ha;
		memory[16'h6ce8] <= 8'ha0;
		memory[16'h6ce9] <= 8'h2e;
		memory[16'h6cea] <= 8'haf;
		memory[16'h6ceb] <= 8'h82;
		memory[16'h6cec] <= 8'h99;
		memory[16'h6ced] <= 8'h99;
		memory[16'h6cee] <= 8'h41;
		memory[16'h6cef] <= 8'h2e;
		memory[16'h6cf0] <= 8'h9c;
		memory[16'h6cf1] <= 8'hb9;
		memory[16'h6cf2] <= 8'hf1;
		memory[16'h6cf3] <= 8'h6c;
		memory[16'h6cf4] <= 8'h3b;
		memory[16'h6cf5] <= 8'hdb;
		memory[16'h6cf6] <= 8'hec;
		memory[16'h6cf7] <= 8'h23;
		memory[16'h6cf8] <= 8'h26;
		memory[16'h6cf9] <= 8'h82;
		memory[16'h6cfa] <= 8'hd8;
		memory[16'h6cfb] <= 8'hc3;
		memory[16'h6cfc] <= 8'h9b;
		memory[16'h6cfd] <= 8'h77;
		memory[16'h6cfe] <= 8'h13;
		memory[16'h6cff] <= 8'h3f;
		memory[16'h6d00] <= 8'h4e;
		memory[16'h6d01] <= 8'ha7;
		memory[16'h6d02] <= 8'h5b;
		memory[16'h6d03] <= 8'h8c;
		memory[16'h6d04] <= 8'h43;
		memory[16'h6d05] <= 8'h2b;
		memory[16'h6d06] <= 8'h96;
		memory[16'h6d07] <= 8'he4;
		memory[16'h6d08] <= 8'h5a;
		memory[16'h6d09] <= 8'h45;
		memory[16'h6d0a] <= 8'h66;
		memory[16'h6d0b] <= 8'hf3;
		memory[16'h6d0c] <= 8'hde;
		memory[16'h6d0d] <= 8'ha8;
		memory[16'h6d0e] <= 8'h21;
		memory[16'h6d0f] <= 8'h7a;
		memory[16'h6d10] <= 8'h61;
		memory[16'h6d11] <= 8'h13;
		memory[16'h6d12] <= 8'he6;
		memory[16'h6d13] <= 8'h9c;
		memory[16'h6d14] <= 8'hee;
		memory[16'h6d15] <= 8'hd3;
		memory[16'h6d16] <= 8'hbf;
		memory[16'h6d17] <= 8'h14;
		memory[16'h6d18] <= 8'h55;
		memory[16'h6d19] <= 8'h97;
		memory[16'h6d1a] <= 8'hd8;
		memory[16'h6d1b] <= 8'hf1;
		memory[16'h6d1c] <= 8'he;
		memory[16'h6d1d] <= 8'heb;
		memory[16'h6d1e] <= 8'h30;
		memory[16'h6d1f] <= 8'h5c;
		memory[16'h6d20] <= 8'h93;
		memory[16'h6d21] <= 8'h8b;
		memory[16'h6d22] <= 8'he9;
		memory[16'h6d23] <= 8'hd6;
		memory[16'h6d24] <= 8'hb7;
		memory[16'h6d25] <= 8'h7f;
		memory[16'h6d26] <= 8'hba;
		memory[16'h6d27] <= 8'h11;
		memory[16'h6d28] <= 8'hc5;
		memory[16'h6d29] <= 8'h21;
		memory[16'h6d2a] <= 8'h4;
		memory[16'h6d2b] <= 8'ha3;
		memory[16'h6d2c] <= 8'hc9;
		memory[16'h6d2d] <= 8'h26;
		memory[16'h6d2e] <= 8'h1e;
		memory[16'h6d2f] <= 8'h2a;
		memory[16'h6d30] <= 8'h39;
		memory[16'h6d31] <= 8'h4;
		memory[16'h6d32] <= 8'hc7;
		memory[16'h6d33] <= 8'h27;
		memory[16'h6d34] <= 8'hd7;
		memory[16'h6d35] <= 8'h86;
		memory[16'h6d36] <= 8'h3c;
		memory[16'h6d37] <= 8'h2d;
		memory[16'h6d38] <= 8'h1e;
		memory[16'h6d39] <= 8'h14;
		memory[16'h6d3a] <= 8'h1e;
		memory[16'h6d3b] <= 8'h2c;
		memory[16'h6d3c] <= 8'hff;
		memory[16'h6d3d] <= 8'h4e;
		memory[16'h6d3e] <= 8'h89;
		memory[16'h6d3f] <= 8'h92;
		memory[16'h6d40] <= 8'hda;
		memory[16'h6d41] <= 8'h72;
		memory[16'h6d42] <= 8'h69;
		memory[16'h6d43] <= 8'h91;
		memory[16'h6d44] <= 8'hf1;
		memory[16'h6d45] <= 8'h23;
		memory[16'h6d46] <= 8'ha2;
		memory[16'h6d47] <= 8'hb6;
		memory[16'h6d48] <= 8'h44;
		memory[16'h6d49] <= 8'ha6;
		memory[16'h6d4a] <= 8'h5a;
		memory[16'h6d4b] <= 8'hd;
		memory[16'h6d4c] <= 8'hcc;
		memory[16'h6d4d] <= 8'h78;
		memory[16'h6d4e] <= 8'h38;
		memory[16'h6d4f] <= 8'h5;
		memory[16'h6d50] <= 8'h7c;
		memory[16'h6d51] <= 8'hff;
		memory[16'h6d52] <= 8'h2d;
		memory[16'h6d53] <= 8'h54;
		memory[16'h6d54] <= 8'h85;
		memory[16'h6d55] <= 8'h69;
		memory[16'h6d56] <= 8'h81;
		memory[16'h6d57] <= 8'ha3;
		memory[16'h6d58] <= 8'h7d;
		memory[16'h6d59] <= 8'h9f;
		memory[16'h6d5a] <= 8'hd0;
		memory[16'h6d5b] <= 8'h7c;
		memory[16'h6d5c] <= 8'hed;
		memory[16'h6d5d] <= 8'h59;
		memory[16'h6d5e] <= 8'hf;
		memory[16'h6d5f] <= 8'hc7;
		memory[16'h6d60] <= 8'hcb;
		memory[16'h6d61] <= 8'h78;
		memory[16'h6d62] <= 8'h58;
		memory[16'h6d63] <= 8'hbc;
		memory[16'h6d64] <= 8'h9b;
		memory[16'h6d65] <= 8'hfa;
		memory[16'h6d66] <= 8'h73;
		memory[16'h6d67] <= 8'he0;
		memory[16'h6d68] <= 8'ha1;
		memory[16'h6d69] <= 8'hcd;
		memory[16'h6d6a] <= 8'hed;
		memory[16'h6d6b] <= 8'h6d;
		memory[16'h6d6c] <= 8'h45;
		memory[16'h6d6d] <= 8'h25;
		memory[16'h6d6e] <= 8'h73;
		memory[16'h6d6f] <= 8'hc1;
		memory[16'h6d70] <= 8'h24;
		memory[16'h6d71] <= 8'ha0;
		memory[16'h6d72] <= 8'h15;
		memory[16'h6d73] <= 8'haa;
		memory[16'h6d74] <= 8'h9;
		memory[16'h6d75] <= 8'h96;
		memory[16'h6d76] <= 8'h4d;
		memory[16'h6d77] <= 8'h86;
		memory[16'h6d78] <= 8'h35;
		memory[16'h6d79] <= 8'h1d;
		memory[16'h6d7a] <= 8'h2;
		memory[16'h6d7b] <= 8'h23;
		memory[16'h6d7c] <= 8'h76;
		memory[16'h6d7d] <= 8'h11;
		memory[16'h6d7e] <= 8'hea;
		memory[16'h6d7f] <= 8'h41;
		memory[16'h6d80] <= 8'h89;
		memory[16'h6d81] <= 8'h43;
		memory[16'h6d82] <= 8'hfe;
		memory[16'h6d83] <= 8'h25;
		memory[16'h6d84] <= 8'h3d;
		memory[16'h6d85] <= 8'h71;
		memory[16'h6d86] <= 8'h5;
		memory[16'h6d87] <= 8'hde;
		memory[16'h6d88] <= 8'h3e;
		memory[16'h6d89] <= 8'hf2;
		memory[16'h6d8a] <= 8'h4c;
		memory[16'h6d8b] <= 8'h83;
		memory[16'h6d8c] <= 8'h18;
		memory[16'h6d8d] <= 8'hbf;
		memory[16'h6d8e] <= 8'h44;
		memory[16'h6d8f] <= 8'h3c;
		memory[16'h6d90] <= 8'h5f;
		memory[16'h6d91] <= 8'h5a;
		memory[16'h6d92] <= 8'he6;
		memory[16'h6d93] <= 8'h68;
		memory[16'h6d94] <= 8'hf0;
		memory[16'h6d95] <= 8'h34;
		memory[16'h6d96] <= 8'hee;
		memory[16'h6d97] <= 8'h26;
		memory[16'h6d98] <= 8'h51;
		memory[16'h6d99] <= 8'hf0;
		memory[16'h6d9a] <= 8'h49;
		memory[16'h6d9b] <= 8'hc8;
		memory[16'h6d9c] <= 8'h2;
		memory[16'h6d9d] <= 8'h33;
		memory[16'h6d9e] <= 8'h9;
		memory[16'h6d9f] <= 8'h8b;
		memory[16'h6da0] <= 8'h76;
		memory[16'h6da1] <= 8'h7;
		memory[16'h6da2] <= 8'hb0;
		memory[16'h6da3] <= 8'hb4;
		memory[16'h6da4] <= 8'h78;
		memory[16'h6da5] <= 8'hb5;
		memory[16'h6da6] <= 8'h92;
		memory[16'h6da7] <= 8'hb6;
		memory[16'h6da8] <= 8'ha8;
		memory[16'h6da9] <= 8'hde;
		memory[16'h6daa] <= 8'h39;
		memory[16'h6dab] <= 8'hc0;
		memory[16'h6dac] <= 8'h9d;
		memory[16'h6dad] <= 8'h7e;
		memory[16'h6dae] <= 8'hfc;
		memory[16'h6daf] <= 8'hfc;
		memory[16'h6db0] <= 8'hd8;
		memory[16'h6db1] <= 8'he3;
		memory[16'h6db2] <= 8'h64;
		memory[16'h6db3] <= 8'hc8;
		memory[16'h6db4] <= 8'h17;
		memory[16'h6db5] <= 8'h52;
		memory[16'h6db6] <= 8'hee;
		memory[16'h6db7] <= 8'h68;
		memory[16'h6db8] <= 8'h43;
		memory[16'h6db9] <= 8'h37;
		memory[16'h6dba] <= 8'h30;
		memory[16'h6dbb] <= 8'h45;
		memory[16'h6dbc] <= 8'h6b;
		memory[16'h6dbd] <= 8'h3a;
		memory[16'h6dbe] <= 8'hd0;
		memory[16'h6dbf] <= 8'he1;
		memory[16'h6dc0] <= 8'h41;
		memory[16'h6dc1] <= 8'h81;
		memory[16'h6dc2] <= 8'h95;
		memory[16'h6dc3] <= 8'hba;
		memory[16'h6dc4] <= 8'h36;
		memory[16'h6dc5] <= 8'h28;
		memory[16'h6dc6] <= 8'h70;
		memory[16'h6dc7] <= 8'hde;
		memory[16'h6dc8] <= 8'h6;
		memory[16'h6dc9] <= 8'haa;
		memory[16'h6dca] <= 8'h9e;
		memory[16'h6dcb] <= 8'ha4;
		memory[16'h6dcc] <= 8'h28;
		memory[16'h6dcd] <= 8'h9b;
		memory[16'h6dce] <= 8'ha0;
		memory[16'h6dcf] <= 8'h0;
		memory[16'h6dd0] <= 8'h7e;
		memory[16'h6dd1] <= 8'h5;
		memory[16'h6dd2] <= 8'hc8;
		memory[16'h6dd3] <= 8'h95;
		memory[16'h6dd4] <= 8'h57;
		memory[16'h6dd5] <= 8'hb7;
		memory[16'h6dd6] <= 8'hfd;
		memory[16'h6dd7] <= 8'h9a;
		memory[16'h6dd8] <= 8'hee;
		memory[16'h6dd9] <= 8'h2e;
		memory[16'h6dda] <= 8'hdf;
		memory[16'h6ddb] <= 8'h59;
		memory[16'h6ddc] <= 8'h68;
		memory[16'h6ddd] <= 8'hb0;
		memory[16'h6dde] <= 8'h3b;
		memory[16'h6ddf] <= 8'ha9;
		memory[16'h6de0] <= 8'h31;
		memory[16'h6de1] <= 8'hd0;
		memory[16'h6de2] <= 8'h63;
		memory[16'h6de3] <= 8'h67;
		memory[16'h6de4] <= 8'hf8;
		memory[16'h6de5] <= 8'hd4;
		memory[16'h6de6] <= 8'h46;
		memory[16'h6de7] <= 8'hff;
		memory[16'h6de8] <= 8'h7e;
		memory[16'h6de9] <= 8'he4;
		memory[16'h6dea] <= 8'ha3;
		memory[16'h6deb] <= 8'ha6;
		memory[16'h6dec] <= 8'h7f;
		memory[16'h6ded] <= 8'h43;
		memory[16'h6dee] <= 8'ha6;
		memory[16'h6def] <= 8'hfd;
		memory[16'h6df0] <= 8'h48;
		memory[16'h6df1] <= 8'h6e;
		memory[16'h6df2] <= 8'h92;
		memory[16'h6df3] <= 8'ha0;
		memory[16'h6df4] <= 8'h25;
		memory[16'h6df5] <= 8'h90;
		memory[16'h6df6] <= 8'h3a;
		memory[16'h6df7] <= 8'h14;
		memory[16'h6df8] <= 8'hbe;
		memory[16'h6df9] <= 8'h1a;
		memory[16'h6dfa] <= 8'h6d;
		memory[16'h6dfb] <= 8'h26;
		memory[16'h6dfc] <= 8'hca;
		memory[16'h6dfd] <= 8'ha8;
		memory[16'h6dfe] <= 8'hcf;
		memory[16'h6dff] <= 8'hfb;
		memory[16'h6e00] <= 8'h79;
		memory[16'h6e01] <= 8'h33;
		memory[16'h6e02] <= 8'h62;
		memory[16'h6e03] <= 8'h71;
		memory[16'h6e04] <= 8'h7;
		memory[16'h6e05] <= 8'ha8;
		memory[16'h6e06] <= 8'h70;
		memory[16'h6e07] <= 8'h85;
		memory[16'h6e08] <= 8'h8d;
		memory[16'h6e09] <= 8'h13;
		memory[16'h6e0a] <= 8'h2b;
		memory[16'h6e0b] <= 8'hc;
		memory[16'h6e0c] <= 8'h57;
		memory[16'h6e0d] <= 8'hd1;
		memory[16'h6e0e] <= 8'ha;
		memory[16'h6e0f] <= 8'h9f;
		memory[16'h6e10] <= 8'h3f;
		memory[16'h6e11] <= 8'h9c;
		memory[16'h6e12] <= 8'h3f;
		memory[16'h6e13] <= 8'h65;
		memory[16'h6e14] <= 8'h2c;
		memory[16'h6e15] <= 8'h7a;
		memory[16'h6e16] <= 8'h79;
		memory[16'h6e17] <= 8'hea;
		memory[16'h6e18] <= 8'h94;
		memory[16'h6e19] <= 8'he6;
		memory[16'h6e1a] <= 8'h10;
		memory[16'h6e1b] <= 8'h5e;
		memory[16'h6e1c] <= 8'h8f;
		memory[16'h6e1d] <= 8'he0;
		memory[16'h6e1e] <= 8'h59;
		memory[16'h6e1f] <= 8'h8;
		memory[16'h6e20] <= 8'h13;
		memory[16'h6e21] <= 8'hbb;
		memory[16'h6e22] <= 8'h79;
		memory[16'h6e23] <= 8'h1a;
		memory[16'h6e24] <= 8'h64;
		memory[16'h6e25] <= 8'hea;
		memory[16'h6e26] <= 8'h9f;
		memory[16'h6e27] <= 8'hf1;
		memory[16'h6e28] <= 8'hfd;
		memory[16'h6e29] <= 8'hca;
		memory[16'h6e2a] <= 8'hfd;
		memory[16'h6e2b] <= 8'h54;
		memory[16'h6e2c] <= 8'h9b;
		memory[16'h6e2d] <= 8'h7;
		memory[16'h6e2e] <= 8'hf4;
		memory[16'h6e2f] <= 8'hda;
		memory[16'h6e30] <= 8'ha4;
		memory[16'h6e31] <= 8'h33;
		memory[16'h6e32] <= 8'h3f;
		memory[16'h6e33] <= 8'hd0;
		memory[16'h6e34] <= 8'had;
		memory[16'h6e35] <= 8'hb8;
		memory[16'h6e36] <= 8'hbb;
		memory[16'h6e37] <= 8'h41;
		memory[16'h6e38] <= 8'h9f;
		memory[16'h6e39] <= 8'hcb;
		memory[16'h6e3a] <= 8'h9f;
		memory[16'h6e3b] <= 8'h2e;
		memory[16'h6e3c] <= 8'hab;
		memory[16'h6e3d] <= 8'hf8;
		memory[16'h6e3e] <= 8'h36;
		memory[16'h6e3f] <= 8'hbe;
		memory[16'h6e40] <= 8'hb4;
		memory[16'h6e41] <= 8'haf;
		memory[16'h6e42] <= 8'hd8;
		memory[16'h6e43] <= 8'h18;
		memory[16'h6e44] <= 8'h99;
		memory[16'h6e45] <= 8'h77;
		memory[16'h6e46] <= 8'h9;
		memory[16'h6e47] <= 8'h97;
		memory[16'h6e48] <= 8'h41;
		memory[16'h6e49] <= 8'h6;
		memory[16'h6e4a] <= 8'heb;
		memory[16'h6e4b] <= 8'hdc;
		memory[16'h6e4c] <= 8'he;
		memory[16'h6e4d] <= 8'hdf;
		memory[16'h6e4e] <= 8'hb7;
		memory[16'h6e4f] <= 8'hb2;
		memory[16'h6e50] <= 8'h13;
		memory[16'h6e51] <= 8'hf6;
		memory[16'h6e52] <= 8'h82;
		memory[16'h6e53] <= 8'hc0;
		memory[16'h6e54] <= 8'haf;
		memory[16'h6e55] <= 8'h3d;
		memory[16'h6e56] <= 8'h2;
		memory[16'h6e57] <= 8'h4e;
		memory[16'h6e58] <= 8'h9;
		memory[16'h6e59] <= 8'ha1;
		memory[16'h6e5a] <= 8'h7c;
		memory[16'h6e5b] <= 8'hb4;
		memory[16'h6e5c] <= 8'h9a;
		memory[16'h6e5d] <= 8'hb2;
		memory[16'h6e5e] <= 8'h73;
		memory[16'h6e5f] <= 8'h4e;
		memory[16'h6e60] <= 8'h61;
		memory[16'h6e61] <= 8'h4b;
		memory[16'h6e62] <= 8'h66;
		memory[16'h6e63] <= 8'hfb;
		memory[16'h6e64] <= 8'hc3;
		memory[16'h6e65] <= 8'h6f;
		memory[16'h6e66] <= 8'h92;
		memory[16'h6e67] <= 8'h4;
		memory[16'h6e68] <= 8'h75;
		memory[16'h6e69] <= 8'h7d;
		memory[16'h6e6a] <= 8'he1;
		memory[16'h6e6b] <= 8'h83;
		memory[16'h6e6c] <= 8'h5d;
		memory[16'h6e6d] <= 8'h98;
		memory[16'h6e6e] <= 8'h35;
		memory[16'h6e6f] <= 8'h70;
		memory[16'h6e70] <= 8'h8e;
		memory[16'h6e71] <= 8'hb8;
		memory[16'h6e72] <= 8'h30;
		memory[16'h6e73] <= 8'h3d;
		memory[16'h6e74] <= 8'hf5;
		memory[16'h6e75] <= 8'h32;
		memory[16'h6e76] <= 8'h8b;
		memory[16'h6e77] <= 8'hfe;
		memory[16'h6e78] <= 8'hd4;
		memory[16'h6e79] <= 8'h7;
		memory[16'h6e7a] <= 8'hb3;
		memory[16'h6e7b] <= 8'h6e;
		memory[16'h6e7c] <= 8'hb9;
		memory[16'h6e7d] <= 8'h26;
		memory[16'h6e7e] <= 8'hbc;
		memory[16'h6e7f] <= 8'h1b;
		memory[16'h6e80] <= 8'h71;
		memory[16'h6e81] <= 8'h22;
		memory[16'h6e82] <= 8'h16;
		memory[16'h6e83] <= 8'h34;
		memory[16'h6e84] <= 8'h91;
		memory[16'h6e85] <= 8'ha8;
		memory[16'h6e86] <= 8'h39;
		memory[16'h6e87] <= 8'h6;
		memory[16'h6e88] <= 8'h25;
		memory[16'h6e89] <= 8'h1a;
		memory[16'h6e8a] <= 8'h8a;
		memory[16'h6e8b] <= 8'h82;
		memory[16'h6e8c] <= 8'hb2;
		memory[16'h6e8d] <= 8'hbf;
		memory[16'h6e8e] <= 8'hf2;
		memory[16'h6e8f] <= 8'h40;
		memory[16'h6e90] <= 8'h77;
		memory[16'h6e91] <= 8'h23;
		memory[16'h6e92] <= 8'h7e;
		memory[16'h6e93] <= 8'h6d;
		memory[16'h6e94] <= 8'h55;
		memory[16'h6e95] <= 8'h9;
		memory[16'h6e96] <= 8'h6b;
		memory[16'h6e97] <= 8'h29;
		memory[16'h6e98] <= 8'h11;
		memory[16'h6e99] <= 8'h1e;
		memory[16'h6e9a] <= 8'h97;
		memory[16'h6e9b] <= 8'hca;
		memory[16'h6e9c] <= 8'h44;
		memory[16'h6e9d] <= 8'h53;
		memory[16'h6e9e] <= 8'he5;
		memory[16'h6e9f] <= 8'hb6;
		memory[16'h6ea0] <= 8'h75;
		memory[16'h6ea1] <= 8'hfb;
		memory[16'h6ea2] <= 8'hea;
		memory[16'h6ea3] <= 8'h6;
		memory[16'h6ea4] <= 8'ha3;
		memory[16'h6ea5] <= 8'h23;
		memory[16'h6ea6] <= 8'hd;
		memory[16'h6ea7] <= 8'hc9;
		memory[16'h6ea8] <= 8'h3d;
		memory[16'h6ea9] <= 8'h97;
		memory[16'h6eaa] <= 8'h4b;
		memory[16'h6eab] <= 8'hef;
		memory[16'h6eac] <= 8'h56;
		memory[16'h6ead] <= 8'h3e;
		memory[16'h6eae] <= 8'h30;
		memory[16'h6eaf] <= 8'hce;
		memory[16'h6eb0] <= 8'h61;
		memory[16'h6eb1] <= 8'hae;
		memory[16'h6eb2] <= 8'h3b;
		memory[16'h6eb3] <= 8'hb6;
		memory[16'h6eb4] <= 8'hb7;
		memory[16'h6eb5] <= 8'ha6;
		memory[16'h6eb6] <= 8'he0;
		memory[16'h6eb7] <= 8'hc8;
		memory[16'h6eb8] <= 8'hc5;
		memory[16'h6eb9] <= 8'h77;
		memory[16'h6eba] <= 8'h93;
		memory[16'h6ebb] <= 8'h9;
		memory[16'h6ebc] <= 8'hcb;
		memory[16'h6ebd] <= 8'h78;
		memory[16'h6ebe] <= 8'hbf;
		memory[16'h6ebf] <= 8'h40;
		memory[16'h6ec0] <= 8'h74;
		memory[16'h6ec1] <= 8'haa;
		memory[16'h6ec2] <= 8'h47;
		memory[16'h6ec3] <= 8'h17;
		memory[16'h6ec4] <= 8'hcd;
		memory[16'h6ec5] <= 8'h54;
		memory[16'h6ec6] <= 8'he0;
		memory[16'h6ec7] <= 8'hb;
		memory[16'h6ec8] <= 8'heb;
		memory[16'h6ec9] <= 8'h2c;
		memory[16'h6eca] <= 8'hfa;
		memory[16'h6ecb] <= 8'h41;
		memory[16'h6ecc] <= 8'h6a;
		memory[16'h6ecd] <= 8'h2a;
		memory[16'h6ece] <= 8'hf;
		memory[16'h6ecf] <= 8'hcb;
		memory[16'h6ed0] <= 8'hd8;
		memory[16'h6ed1] <= 8'h4a;
		memory[16'h6ed2] <= 8'h81;
		memory[16'h6ed3] <= 8'h90;
		memory[16'h6ed4] <= 8'hf1;
		memory[16'h6ed5] <= 8'h61;
		memory[16'h6ed6] <= 8'h58;
		memory[16'h6ed7] <= 8'hb6;
		memory[16'h6ed8] <= 8'hd9;
		memory[16'h6ed9] <= 8'heb;
		memory[16'h6eda] <= 8'hbf;
		memory[16'h6edb] <= 8'ha4;
		memory[16'h6edc] <= 8'h64;
		memory[16'h6edd] <= 8'h7f;
		memory[16'h6ede] <= 8'he4;
		memory[16'h6edf] <= 8'hd8;
		memory[16'h6ee0] <= 8'h29;
		memory[16'h6ee1] <= 8'h2b;
		memory[16'h6ee2] <= 8'hef;
		memory[16'h6ee3] <= 8'hf6;
		memory[16'h6ee4] <= 8'h7f;
		memory[16'h6ee5] <= 8'hd0;
		memory[16'h6ee6] <= 8'h1;
		memory[16'h6ee7] <= 8'h6a;
		memory[16'h6ee8] <= 8'hfc;
		memory[16'h6ee9] <= 8'hfc;
		memory[16'h6eea] <= 8'hac;
		memory[16'h6eeb] <= 8'h66;
		memory[16'h6eec] <= 8'h26;
		memory[16'h6eed] <= 8'hbb;
		memory[16'h6eee] <= 8'h31;
		memory[16'h6eef] <= 8'hff;
		memory[16'h6ef0] <= 8'h6;
		memory[16'h6ef1] <= 8'hb2;
		memory[16'h6ef2] <= 8'h8f;
		memory[16'h6ef3] <= 8'hf7;
		memory[16'h6ef4] <= 8'h14;
		memory[16'h6ef5] <= 8'he7;
		memory[16'h6ef6] <= 8'had;
		memory[16'h6ef7] <= 8'hed;
		memory[16'h6ef8] <= 8'hd3;
		memory[16'h6ef9] <= 8'h6c;
		memory[16'h6efa] <= 8'h91;
		memory[16'h6efb] <= 8'h37;
		memory[16'h6efc] <= 8'heb;
		memory[16'h6efd] <= 8'h75;
		memory[16'h6efe] <= 8'hf;
		memory[16'h6eff] <= 8'h14;
		memory[16'h6f00] <= 8'ha1;
		memory[16'h6f01] <= 8'hfe;
		memory[16'h6f02] <= 8'hb;
		memory[16'h6f03] <= 8'h20;
		memory[16'h6f04] <= 8'hce;
		memory[16'h6f05] <= 8'hc;
		memory[16'h6f06] <= 8'h8b;
		memory[16'h6f07] <= 8'hca;
		memory[16'h6f08] <= 8'h8;
		memory[16'h6f09] <= 8'h37;
		memory[16'h6f0a] <= 8'h30;
		memory[16'h6f0b] <= 8'h2f;
		memory[16'h6f0c] <= 8'hf2;
		memory[16'h6f0d] <= 8'h61;
		memory[16'h6f0e] <= 8'h2e;
		memory[16'h6f0f] <= 8'hf8;
		memory[16'h6f10] <= 8'h14;
		memory[16'h6f11] <= 8'hbd;
		memory[16'h6f12] <= 8'hef;
		memory[16'h6f13] <= 8'h28;
		memory[16'h6f14] <= 8'ha4;
		memory[16'h6f15] <= 8'h9c;
		memory[16'h6f16] <= 8'h15;
		memory[16'h6f17] <= 8'h77;
		memory[16'h6f18] <= 8'h9;
		memory[16'h6f19] <= 8'ha6;
		memory[16'h6f1a] <= 8'hae;
		memory[16'h6f1b] <= 8'hf4;
		memory[16'h6f1c] <= 8'h1b;
		memory[16'h6f1d] <= 8'hbd;
		memory[16'h6f1e] <= 8'h9;
		memory[16'h6f1f] <= 8'hbc;
		memory[16'h6f20] <= 8'hbc;
		memory[16'h6f21] <= 8'h14;
		memory[16'h6f22] <= 8'hdd;
		memory[16'h6f23] <= 8'h8a;
		memory[16'h6f24] <= 8'h20;
		memory[16'h6f25] <= 8'h68;
		memory[16'h6f26] <= 8'h55;
		memory[16'h6f27] <= 8'h29;
		memory[16'h6f28] <= 8'h9f;
		memory[16'h6f29] <= 8'h85;
		memory[16'h6f2a] <= 8'h58;
		memory[16'h6f2b] <= 8'h91;
		memory[16'h6f2c] <= 8'he7;
		memory[16'h6f2d] <= 8'h86;
		memory[16'h6f2e] <= 8'h8a;
		memory[16'h6f2f] <= 8'hfb;
		memory[16'h6f30] <= 8'h43;
		memory[16'h6f31] <= 8'h79;
		memory[16'h6f32] <= 8'h23;
		memory[16'h6f33] <= 8'he7;
		memory[16'h6f34] <= 8'h16;
		memory[16'h6f35] <= 8'h38;
		memory[16'h6f36] <= 8'h5f;
		memory[16'h6f37] <= 8'h1f;
		memory[16'h6f38] <= 8'hde;
		memory[16'h6f39] <= 8'hd;
		memory[16'h6f3a] <= 8'h13;
		memory[16'h6f3b] <= 8'hf9;
		memory[16'h6f3c] <= 8'hcb;
		memory[16'h6f3d] <= 8'h1c;
		memory[16'h6f3e] <= 8'hb6;
		memory[16'h6f3f] <= 8'h87;
		memory[16'h6f40] <= 8'h30;
		memory[16'h6f41] <= 8'h93;
		memory[16'h6f42] <= 8'h11;
		memory[16'h6f43] <= 8'h51;
		memory[16'h6f44] <= 8'hfb;
		memory[16'h6f45] <= 8'h66;
		memory[16'h6f46] <= 8'h7a;
		memory[16'h6f47] <= 8'h9a;
		memory[16'h6f48] <= 8'hec;
		memory[16'h6f49] <= 8'hd2;
		memory[16'h6f4a] <= 8'h2b;
		memory[16'h6f4b] <= 8'hd3;
		memory[16'h6f4c] <= 8'h58;
		memory[16'h6f4d] <= 8'hb5;
		memory[16'h6f4e] <= 8'hce;
		memory[16'h6f4f] <= 8'h9b;
		memory[16'h6f50] <= 8'h2f;
		memory[16'h6f51] <= 8'hf1;
		memory[16'h6f52] <= 8'h82;
		memory[16'h6f53] <= 8'h45;
		memory[16'h6f54] <= 8'h29;
		memory[16'h6f55] <= 8'he1;
		memory[16'h6f56] <= 8'h64;
		memory[16'h6f57] <= 8'h7;
		memory[16'h6f58] <= 8'hef;
		memory[16'h6f59] <= 8'h77;
		memory[16'h6f5a] <= 8'h0;
		memory[16'h6f5b] <= 8'hba;
		memory[16'h6f5c] <= 8'h94;
		memory[16'h6f5d] <= 8'hb6;
		memory[16'h6f5e] <= 8'h41;
		memory[16'h6f5f] <= 8'hc4;
		memory[16'h6f60] <= 8'h49;
		memory[16'h6f61] <= 8'h52;
		memory[16'h6f62] <= 8'h15;
		memory[16'h6f63] <= 8'h44;
		memory[16'h6f64] <= 8'hb9;
		memory[16'h6f65] <= 8'h8f;
		memory[16'h6f66] <= 8'hde;
		memory[16'h6f67] <= 8'ha5;
		memory[16'h6f68] <= 8'h61;
		memory[16'h6f69] <= 8'ha;
		memory[16'h6f6a] <= 8'h78;
		memory[16'h6f6b] <= 8'hb9;
		memory[16'h6f6c] <= 8'hbf;
		memory[16'h6f6d] <= 8'h46;
		memory[16'h6f6e] <= 8'h54;
		memory[16'h6f6f] <= 8'hee;
		memory[16'h6f70] <= 8'h37;
		memory[16'h6f71] <= 8'hd7;
		memory[16'h6f72] <= 8'h33;
		memory[16'h6f73] <= 8'h60;
		memory[16'h6f74] <= 8'hb8;
		memory[16'h6f75] <= 8'h97;
		memory[16'h6f76] <= 8'h67;
		memory[16'h6f77] <= 8'ha7;
		memory[16'h6f78] <= 8'hf;
		memory[16'h6f79] <= 8'h67;
		memory[16'h6f7a] <= 8'h61;
		memory[16'h6f7b] <= 8'ha3;
		memory[16'h6f7c] <= 8'h1e;
		memory[16'h6f7d] <= 8'ha2;
		memory[16'h6f7e] <= 8'h67;
		memory[16'h6f7f] <= 8'h67;
		memory[16'h6f80] <= 8'hf5;
		memory[16'h6f81] <= 8'h7d;
		memory[16'h6f82] <= 8'hac;
		memory[16'h6f83] <= 8'hae;
		memory[16'h6f84] <= 8'hc;
		memory[16'h6f85] <= 8'h8a;
		memory[16'h6f86] <= 8'h53;
		memory[16'h6f87] <= 8'h6e;
		memory[16'h6f88] <= 8'h94;
		memory[16'h6f89] <= 8'hcb;
		memory[16'h6f8a] <= 8'h27;
		memory[16'h6f8b] <= 8'h54;
		memory[16'h6f8c] <= 8'h11;
		memory[16'h6f8d] <= 8'h7c;
		memory[16'h6f8e] <= 8'h42;
		memory[16'h6f8f] <= 8'h48;
		memory[16'h6f90] <= 8'h53;
		memory[16'h6f91] <= 8'h76;
		memory[16'h6f92] <= 8'ha8;
		memory[16'h6f93] <= 8'hb;
		memory[16'h6f94] <= 8'hd;
		memory[16'h6f95] <= 8'hf;
		memory[16'h6f96] <= 8'hb3;
		memory[16'h6f97] <= 8'h1c;
		memory[16'h6f98] <= 8'h76;
		memory[16'h6f99] <= 8'h14;
		memory[16'h6f9a] <= 8'hbf;
		memory[16'h6f9b] <= 8'h94;
		memory[16'h6f9c] <= 8'hb7;
		memory[16'h6f9d] <= 8'h27;
		memory[16'h6f9e] <= 8'hfc;
		memory[16'h6f9f] <= 8'hac;
		memory[16'h6fa0] <= 8'ha4;
		memory[16'h6fa1] <= 8'ha8;
		memory[16'h6fa2] <= 8'h5a;
		memory[16'h6fa3] <= 8'hb0;
		memory[16'h6fa4] <= 8'h32;
		memory[16'h6fa5] <= 8'had;
		memory[16'h6fa6] <= 8'h1e;
		memory[16'h6fa7] <= 8'hc7;
		memory[16'h6fa8] <= 8'h78;
		memory[16'h6fa9] <= 8'h46;
		memory[16'h6faa] <= 8'h1b;
		memory[16'h6fab] <= 8'h89;
		memory[16'h6fac] <= 8'hc2;
		memory[16'h6fad] <= 8'h5d;
		memory[16'h6fae] <= 8'hd1;
		memory[16'h6faf] <= 8'h15;
		memory[16'h6fb0] <= 8'hd3;
		memory[16'h6fb1] <= 8'h79;
		memory[16'h6fb2] <= 8'h20;
		memory[16'h6fb3] <= 8'he1;
		memory[16'h6fb4] <= 8'h88;
		memory[16'h6fb5] <= 8'hd3;
		memory[16'h6fb6] <= 8'hfd;
		memory[16'h6fb7] <= 8'hfe;
		memory[16'h6fb8] <= 8'he8;
		memory[16'h6fb9] <= 8'hbd;
		memory[16'h6fba] <= 8'h93;
		memory[16'h6fbb] <= 8'h9f;
		memory[16'h6fbc] <= 8'he4;
		memory[16'h6fbd] <= 8'h8f;
		memory[16'h6fbe] <= 8'h4b;
		memory[16'h6fbf] <= 8'h88;
		memory[16'h6fc0] <= 8'h37;
		memory[16'h6fc1] <= 8'ha5;
		memory[16'h6fc2] <= 8'h38;
		memory[16'h6fc3] <= 8'h69;
		memory[16'h6fc4] <= 8'h52;
		memory[16'h6fc5] <= 8'h57;
		memory[16'h6fc6] <= 8'h30;
		memory[16'h6fc7] <= 8'hca;
		memory[16'h6fc8] <= 8'h9d;
		memory[16'h6fc9] <= 8'h4b;
		memory[16'h6fca] <= 8'h53;
		memory[16'h6fcb] <= 8'h5f;
		memory[16'h6fcc] <= 8'ha9;
		memory[16'h6fcd] <= 8'h24;
		memory[16'h6fce] <= 8'h74;
		memory[16'h6fcf] <= 8'h7c;
		memory[16'h6fd0] <= 8'h9d;
		memory[16'h6fd1] <= 8'h94;
		memory[16'h6fd2] <= 8'h5d;
		memory[16'h6fd3] <= 8'h25;
		memory[16'h6fd4] <= 8'h68;
		memory[16'h6fd5] <= 8'h5b;
		memory[16'h6fd6] <= 8'h23;
		memory[16'h6fd7] <= 8'h50;
		memory[16'h6fd8] <= 8'h18;
		memory[16'h6fd9] <= 8'hb6;
		memory[16'h6fda] <= 8'hef;
		memory[16'h6fdb] <= 8'hfc;
		memory[16'h6fdc] <= 8'h45;
		memory[16'h6fdd] <= 8'h3a;
		memory[16'h6fde] <= 8'h84;
		memory[16'h6fdf] <= 8'h7c;
		memory[16'h6fe0] <= 8'hdf;
		memory[16'h6fe1] <= 8'hbc;
		memory[16'h6fe2] <= 8'he6;
		memory[16'h6fe3] <= 8'h31;
		memory[16'h6fe4] <= 8'h13;
		memory[16'h6fe5] <= 8'h16;
		memory[16'h6fe6] <= 8'hfb;
		memory[16'h6fe7] <= 8'hb0;
		memory[16'h6fe8] <= 8'h62;
		memory[16'h6fe9] <= 8'h4e;
		memory[16'h6fea] <= 8'hf;
		memory[16'h6feb] <= 8'hb;
		memory[16'h6fec] <= 8'h72;
		memory[16'h6fed] <= 8'h83;
		memory[16'h6fee] <= 8'h87;
		memory[16'h6fef] <= 8'hf;
		memory[16'h6ff0] <= 8'h18;
		memory[16'h6ff1] <= 8'he5;
		memory[16'h6ff2] <= 8'h34;
		memory[16'h6ff3] <= 8'h80;
		memory[16'h6ff4] <= 8'h40;
		memory[16'h6ff5] <= 8'h57;
		memory[16'h6ff6] <= 8'hd0;
		memory[16'h6ff7] <= 8'h58;
		memory[16'h6ff8] <= 8'he;
		memory[16'h6ff9] <= 8'hbf;
		memory[16'h6ffa] <= 8'h54;
		memory[16'h6ffb] <= 8'h53;
		memory[16'h6ffc] <= 8'hf9;
		memory[16'h6ffd] <= 8'hd8;
		memory[16'h6ffe] <= 8'hd0;
		memory[16'h6fff] <= 8'hd8;
		memory[16'h7000] <= 8'h94;
		memory[16'h7001] <= 8'hb6;
		memory[16'h7002] <= 8'h9;
		memory[16'h7003] <= 8'ha8;
		memory[16'h7004] <= 8'hcc;
		memory[16'h7005] <= 8'h4;
		memory[16'h7006] <= 8'h58;
		memory[16'h7007] <= 8'h2e;
		memory[16'h7008] <= 8'h52;
		memory[16'h7009] <= 8'h68;
		memory[16'h700a] <= 8'h39;
		memory[16'h700b] <= 8'hc4;
		memory[16'h700c] <= 8'heb;
		memory[16'h700d] <= 8'hc1;
		memory[16'h700e] <= 8'hd3;
		memory[16'h700f] <= 8'h3;
		memory[16'h7010] <= 8'ha6;
		memory[16'h7011] <= 8'h7;
		memory[16'h7012] <= 8'h83;
		memory[16'h7013] <= 8'he6;
		memory[16'h7014] <= 8'h5e;
		memory[16'h7015] <= 8'h53;
		memory[16'h7016] <= 8'h3e;
		memory[16'h7017] <= 8'h6c;
		memory[16'h7018] <= 8'h12;
		memory[16'h7019] <= 8'h92;
		memory[16'h701a] <= 8'hc0;
		memory[16'h701b] <= 8'hb;
		memory[16'h701c] <= 8'h6a;
		memory[16'h701d] <= 8'h90;
		memory[16'h701e] <= 8'he3;
		memory[16'h701f] <= 8'hfe;
		memory[16'h7020] <= 8'h46;
		memory[16'h7021] <= 8'hec;
		memory[16'h7022] <= 8'ha6;
		memory[16'h7023] <= 8'h12;
		memory[16'h7024] <= 8'hf0;
		memory[16'h7025] <= 8'hff;
		memory[16'h7026] <= 8'h41;
		memory[16'h7027] <= 8'h42;
		memory[16'h7028] <= 8'h67;
		memory[16'h7029] <= 8'h7a;
		memory[16'h702a] <= 8'h6;
		memory[16'h702b] <= 8'h52;
		memory[16'h702c] <= 8'h3b;
		memory[16'h702d] <= 8'hd9;
		memory[16'h702e] <= 8'h56;
		memory[16'h702f] <= 8'he1;
		memory[16'h7030] <= 8'he0;
		memory[16'h7031] <= 8'hd9;
		memory[16'h7032] <= 8'hc7;
		memory[16'h7033] <= 8'h3f;
		memory[16'h7034] <= 8'h2d;
		memory[16'h7035] <= 8'h5;
		memory[16'h7036] <= 8'hab;
		memory[16'h7037] <= 8'h3f;
		memory[16'h7038] <= 8'h97;
		memory[16'h7039] <= 8'h6b;
		memory[16'h703a] <= 8'h4b;
		memory[16'h703b] <= 8'h1;
		memory[16'h703c] <= 8'hfb;
		memory[16'h703d] <= 8'h2e;
		memory[16'h703e] <= 8'h0;
		memory[16'h703f] <= 8'h41;
		memory[16'h7040] <= 8'h1b;
		memory[16'h7041] <= 8'ha6;
		memory[16'h7042] <= 8'h54;
		memory[16'h7043] <= 8'hb;
		memory[16'h7044] <= 8'ha5;
		memory[16'h7045] <= 8'h95;
		memory[16'h7046] <= 8'h4e;
		memory[16'h7047] <= 8'hc;
		memory[16'h7048] <= 8'hf;
		memory[16'h7049] <= 8'h54;
		memory[16'h704a] <= 8'h5f;
		memory[16'h704b] <= 8'h4b;
		memory[16'h704c] <= 8'h2e;
		memory[16'h704d] <= 8'hb5;
		memory[16'h704e] <= 8'h2c;
		memory[16'h704f] <= 8'he;
		memory[16'h7050] <= 8'h8e;
		memory[16'h7051] <= 8'hf4;
		memory[16'h7052] <= 8'h4d;
		memory[16'h7053] <= 8'hbb;
		memory[16'h7054] <= 8'hf9;
		memory[16'h7055] <= 8'hf9;
		memory[16'h7056] <= 8'hfb;
		memory[16'h7057] <= 8'h91;
		memory[16'h7058] <= 8'h64;
		memory[16'h7059] <= 8'h46;
		memory[16'h705a] <= 8'h92;
		memory[16'h705b] <= 8'h60;
		memory[16'h705c] <= 8'h74;
		memory[16'h705d] <= 8'h92;
		memory[16'h705e] <= 8'ha1;
		memory[16'h705f] <= 8'h8f;
		memory[16'h7060] <= 8'h39;
		memory[16'h7061] <= 8'hf5;
		memory[16'h7062] <= 8'h9b;
		memory[16'h7063] <= 8'hde;
		memory[16'h7064] <= 8'h8a;
		memory[16'h7065] <= 8'he9;
		memory[16'h7066] <= 8'heb;
		memory[16'h7067] <= 8'h9a;
		memory[16'h7068] <= 8'h3d;
		memory[16'h7069] <= 8'h4a;
		memory[16'h706a] <= 8'he5;
		memory[16'h706b] <= 8'h6b;
		memory[16'h706c] <= 8'hff;
		memory[16'h706d] <= 8'h11;
		memory[16'h706e] <= 8'h7a;
		memory[16'h706f] <= 8'h8d;
		memory[16'h7070] <= 8'h5;
		memory[16'h7071] <= 8'hc7;
		memory[16'h7072] <= 8'h49;
		memory[16'h7073] <= 8'hff;
		memory[16'h7074] <= 8'hc0;
		memory[16'h7075] <= 8'h44;
		memory[16'h7076] <= 8'h90;
		memory[16'h7077] <= 8'h25;
		memory[16'h7078] <= 8'h8a;
		memory[16'h7079] <= 8'h22;
		memory[16'h707a] <= 8'h85;
		memory[16'h707b] <= 8'hfe;
		memory[16'h707c] <= 8'hb5;
		memory[16'h707d] <= 8'h26;
		memory[16'h707e] <= 8'h8e;
		memory[16'h707f] <= 8'hee;
		memory[16'h7080] <= 8'h1c;
		memory[16'h7081] <= 8'h29;
		memory[16'h7082] <= 8'hcc;
		memory[16'h7083] <= 8'ha6;
		memory[16'h7084] <= 8'h12;
		memory[16'h7085] <= 8'hb7;
		memory[16'h7086] <= 8'h40;
		memory[16'h7087] <= 8'h4f;
		memory[16'h7088] <= 8'h1;
		memory[16'h7089] <= 8'h25;
		memory[16'h708a] <= 8'hbb;
		memory[16'h708b] <= 8'h0;
		memory[16'h708c] <= 8'h37;
		memory[16'h708d] <= 8'h35;
		memory[16'h708e] <= 8'h8e;
		memory[16'h708f] <= 8'h3c;
		memory[16'h7090] <= 8'hfc;
		memory[16'h7091] <= 8'hd7;
		memory[16'h7092] <= 8'h3b;
		memory[16'h7093] <= 8'hbd;
		memory[16'h7094] <= 8'h1b;
		memory[16'h7095] <= 8'hcb;
		memory[16'h7096] <= 8'he2;
		memory[16'h7097] <= 8'ha5;
		memory[16'h7098] <= 8'hee;
		memory[16'h7099] <= 8'h67;
		memory[16'h709a] <= 8'ha3;
		memory[16'h709b] <= 8'ha3;
		memory[16'h709c] <= 8'h8d;
		memory[16'h709d] <= 8'h31;
		memory[16'h709e] <= 8'h91;
		memory[16'h709f] <= 8'ha9;
		memory[16'h70a0] <= 8'h5a;
		memory[16'h70a1] <= 8'h5d;
		memory[16'h70a2] <= 8'h50;
		memory[16'h70a3] <= 8'h6c;
		memory[16'h70a4] <= 8'h15;
		memory[16'h70a5] <= 8'h90;
		memory[16'h70a6] <= 8'hbc;
		memory[16'h70a7] <= 8'h16;
		memory[16'h70a8] <= 8'hb6;
		memory[16'h70a9] <= 8'h77;
		memory[16'h70aa] <= 8'h17;
		memory[16'h70ab] <= 8'hed;
		memory[16'h70ac] <= 8'hac;
		memory[16'h70ad] <= 8'ha5;
		memory[16'h70ae] <= 8'h29;
		memory[16'h70af] <= 8'ha8;
		memory[16'h70b0] <= 8'h7c;
		memory[16'h70b1] <= 8'h65;
		memory[16'h70b2] <= 8'h65;
		memory[16'h70b3] <= 8'h97;
		memory[16'h70b4] <= 8'h30;
		memory[16'h70b5] <= 8'h47;
		memory[16'h70b6] <= 8'h3c;
		memory[16'h70b7] <= 8'h1e;
		memory[16'h70b8] <= 8'hae;
		memory[16'h70b9] <= 8'hdf;
		memory[16'h70ba] <= 8'hc1;
		memory[16'h70bb] <= 8'h3c;
		memory[16'h70bc] <= 8'h11;
		memory[16'h70bd] <= 8'h52;
		memory[16'h70be] <= 8'he5;
		memory[16'h70bf] <= 8'h6b;
		memory[16'h70c0] <= 8'hb0;
		memory[16'h70c1] <= 8'h35;
		memory[16'h70c2] <= 8'hd8;
		memory[16'h70c3] <= 8'hc5;
		memory[16'h70c4] <= 8'hc6;
		memory[16'h70c5] <= 8'h94;
		memory[16'h70c6] <= 8'hdb;
		memory[16'h70c7] <= 8'h7c;
		memory[16'h70c8] <= 8'hb;
		memory[16'h70c9] <= 8'hf2;
		memory[16'h70ca] <= 8'h69;
		memory[16'h70cb] <= 8'hb7;
		memory[16'h70cc] <= 8'h97;
		memory[16'h70cd] <= 8'h92;
		memory[16'h70ce] <= 8'h5f;
		memory[16'h70cf] <= 8'h13;
		memory[16'h70d0] <= 8'hf7;
		memory[16'h70d1] <= 8'hc5;
		memory[16'h70d2] <= 8'haa;
		memory[16'h70d3] <= 8'h28;
		memory[16'h70d4] <= 8'hc;
		memory[16'h70d5] <= 8'he6;
		memory[16'h70d6] <= 8'h46;
		memory[16'h70d7] <= 8'hbb;
		memory[16'h70d8] <= 8'hc6;
		memory[16'h70d9] <= 8'h8;
		memory[16'h70da] <= 8'hf7;
		memory[16'h70db] <= 8'hd7;
		memory[16'h70dc] <= 8'h5a;
		memory[16'h70dd] <= 8'hdc;
		memory[16'h70de] <= 8'h42;
		memory[16'h70df] <= 8'ha;
		memory[16'h70e0] <= 8'h12;
		memory[16'h70e1] <= 8'h1a;
		memory[16'h70e2] <= 8'hcf;
		memory[16'h70e3] <= 8'hd8;
		memory[16'h70e4] <= 8'hae;
		memory[16'h70e5] <= 8'hab;
		memory[16'h70e6] <= 8'h54;
		memory[16'h70e7] <= 8'hb9;
		memory[16'h70e8] <= 8'h9d;
		memory[16'h70e9] <= 8'hbd;
		memory[16'h70ea] <= 8'h70;
		memory[16'h70eb] <= 8'h35;
		memory[16'h70ec] <= 8'h4f;
		memory[16'h70ed] <= 8'hd0;
		memory[16'h70ee] <= 8'h48;
		memory[16'h70ef] <= 8'h47;
		memory[16'h70f0] <= 8'h95;
		memory[16'h70f1] <= 8'hf3;
		memory[16'h70f2] <= 8'h6f;
		memory[16'h70f3] <= 8'ha1;
		memory[16'h70f4] <= 8'hd9;
		memory[16'h70f5] <= 8'hb5;
		memory[16'h70f6] <= 8'h5c;
		memory[16'h70f7] <= 8'h9f;
		memory[16'h70f8] <= 8'hbd;
		memory[16'h70f9] <= 8'h53;
		memory[16'h70fa] <= 8'h76;
		memory[16'h70fb] <= 8'h18;
		memory[16'h70fc] <= 8'h30;
		memory[16'h70fd] <= 8'hb9;
		memory[16'h70fe] <= 8'h22;
		memory[16'h70ff] <= 8'h42;
		memory[16'h7100] <= 8'hd3;
		memory[16'h7101] <= 8'hf2;
		memory[16'h7102] <= 8'h1a;
		memory[16'h7103] <= 8'h82;
		memory[16'h7104] <= 8'h9d;
		memory[16'h7105] <= 8'h6e;
		memory[16'h7106] <= 8'h3b;
		memory[16'h7107] <= 8'h3a;
		memory[16'h7108] <= 8'h2b;
		memory[16'h7109] <= 8'hac;
		memory[16'h710a] <= 8'h6f;
		memory[16'h710b] <= 8'h7a;
		memory[16'h710c] <= 8'h7c;
		memory[16'h710d] <= 8'hb8;
		memory[16'h710e] <= 8'hc1;
		memory[16'h710f] <= 8'h11;
		memory[16'h7110] <= 8'hab;
		memory[16'h7111] <= 8'h30;
		memory[16'h7112] <= 8'hb2;
		memory[16'h7113] <= 8'h84;
		memory[16'h7114] <= 8'he6;
		memory[16'h7115] <= 8'hf;
		memory[16'h7116] <= 8'h24;
		memory[16'h7117] <= 8'ha3;
		memory[16'h7118] <= 8'h62;
		memory[16'h7119] <= 8'h9a;
		memory[16'h711a] <= 8'hbb;
		memory[16'h711b] <= 8'h92;
		memory[16'h711c] <= 8'h53;
		memory[16'h711d] <= 8'hde;
		memory[16'h711e] <= 8'hd4;
		memory[16'h711f] <= 8'h27;
		memory[16'h7120] <= 8'hd0;
		memory[16'h7121] <= 8'hee;
		memory[16'h7122] <= 8'ha9;
		memory[16'h7123] <= 8'h6d;
		memory[16'h7124] <= 8'h5c;
		memory[16'h7125] <= 8'he4;
		memory[16'h7126] <= 8'ha7;
		memory[16'h7127] <= 8'h87;
		memory[16'h7128] <= 8'h90;
		memory[16'h7129] <= 8'h17;
		memory[16'h712a] <= 8'h2;
		memory[16'h712b] <= 8'hc;
		memory[16'h712c] <= 8'hcf;
		memory[16'h712d] <= 8'hc3;
		memory[16'h712e] <= 8'h1d;
		memory[16'h712f] <= 8'h7a;
		memory[16'h7130] <= 8'hf4;
		memory[16'h7131] <= 8'hd0;
		memory[16'h7132] <= 8'hfe;
		memory[16'h7133] <= 8'hda;
		memory[16'h7134] <= 8'hdf;
		memory[16'h7135] <= 8'h22;
		memory[16'h7136] <= 8'h7d;
		memory[16'h7137] <= 8'h41;
		memory[16'h7138] <= 8'hbd;
		memory[16'h7139] <= 8'h39;
		memory[16'h713a] <= 8'hd4;
		memory[16'h713b] <= 8'h10;
		memory[16'h713c] <= 8'h17;
		memory[16'h713d] <= 8'ha8;
		memory[16'h713e] <= 8'h37;
		memory[16'h713f] <= 8'he7;
		memory[16'h7140] <= 8'h97;
		memory[16'h7141] <= 8'he0;
		memory[16'h7142] <= 8'h54;
		memory[16'h7143] <= 8'hf3;
		memory[16'h7144] <= 8'hc5;
		memory[16'h7145] <= 8'hfb;
		memory[16'h7146] <= 8'h7b;
		memory[16'h7147] <= 8'h55;
		memory[16'h7148] <= 8'h12;
		memory[16'h7149] <= 8'h7d;
		memory[16'h714a] <= 8'h62;
		memory[16'h714b] <= 8'he1;
		memory[16'h714c] <= 8'h40;
		memory[16'h714d] <= 8'h7f;
		memory[16'h714e] <= 8'h5b;
		memory[16'h714f] <= 8'h34;
		memory[16'h7150] <= 8'h4f;
		memory[16'h7151] <= 8'h5a;
		memory[16'h7152] <= 8'he;
		memory[16'h7153] <= 8'h2e;
		memory[16'h7154] <= 8'h7c;
		memory[16'h7155] <= 8'h8c;
		memory[16'h7156] <= 8'h70;
		memory[16'h7157] <= 8'h39;
		memory[16'h7158] <= 8'hc5;
		memory[16'h7159] <= 8'h44;
		memory[16'h715a] <= 8'h4a;
		memory[16'h715b] <= 8'hdc;
		memory[16'h715c] <= 8'hec;
		memory[16'h715d] <= 8'h81;
		memory[16'h715e] <= 8'hc3;
		memory[16'h715f] <= 8'h83;
		memory[16'h7160] <= 8'h62;
		memory[16'h7161] <= 8'h17;
		memory[16'h7162] <= 8'h77;
		memory[16'h7163] <= 8'h27;
		memory[16'h7164] <= 8'h12;
		memory[16'h7165] <= 8'hf2;
		memory[16'h7166] <= 8'h7c;
		memory[16'h7167] <= 8'h25;
		memory[16'h7168] <= 8'h6f;
		memory[16'h7169] <= 8'hde;
		memory[16'h716a] <= 8'h6;
		memory[16'h716b] <= 8'haf;
		memory[16'h716c] <= 8'h5e;
		memory[16'h716d] <= 8'h62;
		memory[16'h716e] <= 8'he4;
		memory[16'h716f] <= 8'had;
		memory[16'h7170] <= 8'hbc;
		memory[16'h7171] <= 8'hf2;
		memory[16'h7172] <= 8'hdc;
		memory[16'h7173] <= 8'h38;
		memory[16'h7174] <= 8'h7e;
		memory[16'h7175] <= 8'h4c;
		memory[16'h7176] <= 8'h72;
		memory[16'h7177] <= 8'h43;
		memory[16'h7178] <= 8'h90;
		memory[16'h7179] <= 8'hbc;
		memory[16'h717a] <= 8'h1f;
		memory[16'h717b] <= 8'h7c;
		memory[16'h717c] <= 8'h3d;
		memory[16'h717d] <= 8'he2;
		memory[16'h717e] <= 8'h0;
		memory[16'h717f] <= 8'h9f;
		memory[16'h7180] <= 8'hf9;
		memory[16'h7181] <= 8'h77;
		memory[16'h7182] <= 8'hc6;
		memory[16'h7183] <= 8'hc;
		memory[16'h7184] <= 8'h69;
		memory[16'h7185] <= 8'h43;
		memory[16'h7186] <= 8'h31;
		memory[16'h7187] <= 8'hd8;
		memory[16'h7188] <= 8'h21;
		memory[16'h7189] <= 8'h37;
		memory[16'h718a] <= 8'h87;
		memory[16'h718b] <= 8'h7f;
		memory[16'h718c] <= 8'h99;
		memory[16'h718d] <= 8'h6b;
		memory[16'h718e] <= 8'h2d;
		memory[16'h718f] <= 8'h55;
		memory[16'h7190] <= 8'h5e;
		memory[16'h7191] <= 8'h9;
		memory[16'h7192] <= 8'h8e;
		memory[16'h7193] <= 8'hdc;
		memory[16'h7194] <= 8'h55;
		memory[16'h7195] <= 8'h0;
		memory[16'h7196] <= 8'h20;
		memory[16'h7197] <= 8'he5;
		memory[16'h7198] <= 8'hbc;
		memory[16'h7199] <= 8'h3f;
		memory[16'h719a] <= 8'h61;
		memory[16'h719b] <= 8'hf9;
		memory[16'h719c] <= 8'h22;
		memory[16'h719d] <= 8'h61;
		memory[16'h719e] <= 8'h99;
		memory[16'h719f] <= 8'h1b;
		memory[16'h71a0] <= 8'hd8;
		memory[16'h71a1] <= 8'h5f;
		memory[16'h71a2] <= 8'h27;
		memory[16'h71a3] <= 8'h41;
		memory[16'h71a4] <= 8'ha2;
		memory[16'h71a5] <= 8'h58;
		memory[16'h71a6] <= 8'h19;
		memory[16'h71a7] <= 8'hc4;
		memory[16'h71a8] <= 8'h90;
		memory[16'h71a9] <= 8'ha1;
		memory[16'h71aa] <= 8'h43;
		memory[16'h71ab] <= 8'h29;
		memory[16'h71ac] <= 8'hc;
		memory[16'h71ad] <= 8'h70;
		memory[16'h71ae] <= 8'h7f;
		memory[16'h71af] <= 8'h6a;
		memory[16'h71b0] <= 8'h79;
		memory[16'h71b1] <= 8'hd;
		memory[16'h71b2] <= 8'h47;
		memory[16'h71b3] <= 8'hce;
		memory[16'h71b4] <= 8'hd;
		memory[16'h71b5] <= 8'h67;
		memory[16'h71b6] <= 8'hb3;
		memory[16'h71b7] <= 8'hc9;
		memory[16'h71b8] <= 8'ha6;
		memory[16'h71b9] <= 8'h15;
		memory[16'h71ba] <= 8'hc2;
		memory[16'h71bb] <= 8'hc8;
		memory[16'h71bc] <= 8'h76;
		memory[16'h71bd] <= 8'h5b;
		memory[16'h71be] <= 8'he4;
		memory[16'h71bf] <= 8'h4f;
		memory[16'h71c0] <= 8'hbb;
		memory[16'h71c1] <= 8'hb;
		memory[16'h71c2] <= 8'h90;
		memory[16'h71c3] <= 8'h5d;
		memory[16'h71c4] <= 8'h64;
		memory[16'h71c5] <= 8'haa;
		memory[16'h71c6] <= 8'h21;
		memory[16'h71c7] <= 8'hf4;
		memory[16'h71c8] <= 8'h4b;
		memory[16'h71c9] <= 8'h65;
		memory[16'h71ca] <= 8'h1d;
		memory[16'h71cb] <= 8'h57;
		memory[16'h71cc] <= 8'hd5;
		memory[16'h71cd] <= 8'h9c;
		memory[16'h71ce] <= 8'hc2;
		memory[16'h71cf] <= 8'h4f;
		memory[16'h71d0] <= 8'ha9;
		memory[16'h71d1] <= 8'h9;
		memory[16'h71d2] <= 8'h1d;
		memory[16'h71d3] <= 8'hb6;
		memory[16'h71d4] <= 8'h70;
		memory[16'h71d5] <= 8'hd1;
		memory[16'h71d6] <= 8'h7f;
		memory[16'h71d7] <= 8'h16;
		memory[16'h71d8] <= 8'he6;
		memory[16'h71d9] <= 8'h42;
		memory[16'h71da] <= 8'hdf;
		memory[16'h71db] <= 8'h5c;
		memory[16'h71dc] <= 8'h9d;
		memory[16'h71dd] <= 8'hc3;
		memory[16'h71de] <= 8'hab;
		memory[16'h71df] <= 8'h58;
		memory[16'h71e0] <= 8'hce;
		memory[16'h71e1] <= 8'h3c;
		memory[16'h71e2] <= 8'hb6;
		memory[16'h71e3] <= 8'h32;
		memory[16'h71e4] <= 8'he6;
		memory[16'h71e5] <= 8'hd7;
		memory[16'h71e6] <= 8'h26;
		memory[16'h71e7] <= 8'h31;
		memory[16'h71e8] <= 8'h3c;
		memory[16'h71e9] <= 8'h44;
		memory[16'h71ea] <= 8'h88;
		memory[16'h71eb] <= 8'h12;
		memory[16'h71ec] <= 8'he0;
		memory[16'h71ed] <= 8'h4a;
		memory[16'h71ee] <= 8'h61;
		memory[16'h71ef] <= 8'h8a;
		memory[16'h71f0] <= 8'h53;
		memory[16'h71f1] <= 8'h7e;
		memory[16'h71f2] <= 8'h40;
		memory[16'h71f3] <= 8'hc3;
		memory[16'h71f4] <= 8'h4f;
		memory[16'h71f5] <= 8'hc0;
		memory[16'h71f6] <= 8'hda;
		memory[16'h71f7] <= 8'h35;
		memory[16'h71f8] <= 8'h2;
		memory[16'h71f9] <= 8'hb9;
		memory[16'h71fa] <= 8'h92;
		memory[16'h71fb] <= 8'h9f;
		memory[16'h71fc] <= 8'h7c;
		memory[16'h71fd] <= 8'h3d;
		memory[16'h71fe] <= 8'hf8;
		memory[16'h71ff] <= 8'h4a;
		memory[16'h7200] <= 8'h79;
		memory[16'h7201] <= 8'hae;
		memory[16'h7202] <= 8'h7d;
		memory[16'h7203] <= 8'h5f;
		memory[16'h7204] <= 8'h85;
		memory[16'h7205] <= 8'ha3;
		memory[16'h7206] <= 8'h90;
		memory[16'h7207] <= 8'hc2;
		memory[16'h7208] <= 8'he7;
		memory[16'h7209] <= 8'h19;
		memory[16'h720a] <= 8'hd4;
		memory[16'h720b] <= 8'hc8;
		memory[16'h720c] <= 8'h63;
		memory[16'h720d] <= 8'h35;
		memory[16'h720e] <= 8'h52;
		memory[16'h720f] <= 8'hb7;
		memory[16'h7210] <= 8'hb3;
		memory[16'h7211] <= 8'h92;
		memory[16'h7212] <= 8'h7a;
		memory[16'h7213] <= 8'h3;
		memory[16'h7214] <= 8'h52;
		memory[16'h7215] <= 8'h54;
		memory[16'h7216] <= 8'h38;
		memory[16'h7217] <= 8'h54;
		memory[16'h7218] <= 8'hd;
		memory[16'h7219] <= 8'hca;
		memory[16'h721a] <= 8'hf4;
		memory[16'h721b] <= 8'h89;
		memory[16'h721c] <= 8'h8;
		memory[16'h721d] <= 8'hec;
		memory[16'h721e] <= 8'hd4;
		memory[16'h721f] <= 8'h81;
		memory[16'h7220] <= 8'h9a;
		memory[16'h7221] <= 8'h51;
		memory[16'h7222] <= 8'he1;
		memory[16'h7223] <= 8'h1f;
		memory[16'h7224] <= 8'hf4;
		memory[16'h7225] <= 8'h71;
		memory[16'h7226] <= 8'he1;
		memory[16'h7227] <= 8'hdc;
		memory[16'h7228] <= 8'h8a;
		memory[16'h7229] <= 8'hb5;
		memory[16'h722a] <= 8'ha4;
		memory[16'h722b] <= 8'hee;
		memory[16'h722c] <= 8'hea;
		memory[16'h722d] <= 8'hf6;
		memory[16'h722e] <= 8'ha5;
		memory[16'h722f] <= 8'h9e;
		memory[16'h7230] <= 8'h88;
		memory[16'h7231] <= 8'h1f;
		memory[16'h7232] <= 8'ha1;
		memory[16'h7233] <= 8'hdb;
		memory[16'h7234] <= 8'h74;
		memory[16'h7235] <= 8'hd9;
		memory[16'h7236] <= 8'h2f;
		memory[16'h7237] <= 8'h81;
		memory[16'h7238] <= 8'ha4;
		memory[16'h7239] <= 8'h23;
		memory[16'h723a] <= 8'hb;
		memory[16'h723b] <= 8'hac;
		memory[16'h723c] <= 8'hf;
		memory[16'h723d] <= 8'hdf;
		memory[16'h723e] <= 8'h2d;
		memory[16'h723f] <= 8'ha9;
		memory[16'h7240] <= 8'h30;
		memory[16'h7241] <= 8'he;
		memory[16'h7242] <= 8'hc9;
		memory[16'h7243] <= 8'h24;
		memory[16'h7244] <= 8'h80;
		memory[16'h7245] <= 8'haa;
		memory[16'h7246] <= 8'h0;
		memory[16'h7247] <= 8'ha;
		memory[16'h7248] <= 8'h60;
		memory[16'h7249] <= 8'ha4;
		memory[16'h724a] <= 8'hf8;
		memory[16'h724b] <= 8'h4a;
		memory[16'h724c] <= 8'h9a;
		memory[16'h724d] <= 8'h9d;
		memory[16'h724e] <= 8'he8;
		memory[16'h724f] <= 8'h23;
		memory[16'h7250] <= 8'hbd;
		memory[16'h7251] <= 8'h89;
		memory[16'h7252] <= 8'hfe;
		memory[16'h7253] <= 8'h31;
		memory[16'h7254] <= 8'h63;
		memory[16'h7255] <= 8'h2d;
		memory[16'h7256] <= 8'hb2;
		memory[16'h7257] <= 8'h7;
		memory[16'h7258] <= 8'h51;
		memory[16'h7259] <= 8'hbd;
		memory[16'h725a] <= 8'hb3;
		memory[16'h725b] <= 8'h60;
		memory[16'h725c] <= 8'h9c;
		memory[16'h725d] <= 8'he0;
		memory[16'h725e] <= 8'ha;
		memory[16'h725f] <= 8'hcc;
		memory[16'h7260] <= 8'hef;
		memory[16'h7261] <= 8'hd3;
		memory[16'h7262] <= 8'hf1;
		memory[16'h7263] <= 8'h6f;
		memory[16'h7264] <= 8'h7d;
		memory[16'h7265] <= 8'hf1;
		memory[16'h7266] <= 8'h79;
		memory[16'h7267] <= 8'hdd;
		memory[16'h7268] <= 8'h96;
		memory[16'h7269] <= 8'h72;
		memory[16'h726a] <= 8'h28;
		memory[16'h726b] <= 8'h30;
		memory[16'h726c] <= 8'hf;
		memory[16'h726d] <= 8'h10;
		memory[16'h726e] <= 8'h53;
		memory[16'h726f] <= 8'hcc;
		memory[16'h7270] <= 8'h9a;
		memory[16'h7271] <= 8'h51;
		memory[16'h7272] <= 8'hfd;
		memory[16'h7273] <= 8'hfd;
		memory[16'h7274] <= 8'h7f;
		memory[16'h7275] <= 8'hb0;
		memory[16'h7276] <= 8'h4;
		memory[16'h7277] <= 8'hd0;
		memory[16'h7278] <= 8'h6d;
		memory[16'h7279] <= 8'hb7;
		memory[16'h727a] <= 8'h30;
		memory[16'h727b] <= 8'ha;
		memory[16'h727c] <= 8'h97;
		memory[16'h727d] <= 8'h3a;
		memory[16'h727e] <= 8'hd6;
		memory[16'h727f] <= 8'h86;
		memory[16'h7280] <= 8'hd;
		memory[16'h7281] <= 8'hc7;
		memory[16'h7282] <= 8'hf5;
		memory[16'h7283] <= 8'h8b;
		memory[16'h7284] <= 8'hb9;
		memory[16'h7285] <= 8'h6f;
		memory[16'h7286] <= 8'h68;
		memory[16'h7287] <= 8'h4f;
		memory[16'h7288] <= 8'he1;
		memory[16'h7289] <= 8'h90;
		memory[16'h728a] <= 8'h7f;
		memory[16'h728b] <= 8'hf0;
		memory[16'h728c] <= 8'ha1;
		memory[16'h728d] <= 8'hd3;
		memory[16'h728e] <= 8'hbd;
		memory[16'h728f] <= 8'h3b;
		memory[16'h7290] <= 8'h24;
		memory[16'h7291] <= 8'hba;
		memory[16'h7292] <= 8'h38;
		memory[16'h7293] <= 8'ha3;
		memory[16'h7294] <= 8'h6a;
		memory[16'h7295] <= 8'h3c;
		memory[16'h7296] <= 8'h73;
		memory[16'h7297] <= 8'hd8;
		memory[16'h7298] <= 8'hf3;
		memory[16'h7299] <= 8'ha4;
		memory[16'h729a] <= 8'he2;
		memory[16'h729b] <= 8'h8a;
		memory[16'h729c] <= 8'hde;
		memory[16'h729d] <= 8'hb8;
		memory[16'h729e] <= 8'h11;
		memory[16'h729f] <= 8'hec;
		memory[16'h72a0] <= 8'h80;
		memory[16'h72a1] <= 8'h6;
		memory[16'h72a2] <= 8'h77;
		memory[16'h72a3] <= 8'h39;
		memory[16'h72a4] <= 8'h75;
		memory[16'h72a5] <= 8'hdf;
		memory[16'h72a6] <= 8'h88;
		memory[16'h72a7] <= 8'h56;
		memory[16'h72a8] <= 8'h70;
		memory[16'h72a9] <= 8'h7;
		memory[16'h72aa] <= 8'h47;
		memory[16'h72ab] <= 8'h11;
		memory[16'h72ac] <= 8'hda;
		memory[16'h72ad] <= 8'h4;
		memory[16'h72ae] <= 8'h4c;
		memory[16'h72af] <= 8'hff;
		memory[16'h72b0] <= 8'hbe;
		memory[16'h72b1] <= 8'h84;
		memory[16'h72b2] <= 8'ha2;
		memory[16'h72b3] <= 8'h29;
		memory[16'h72b4] <= 8'hc0;
		memory[16'h72b5] <= 8'h16;
		memory[16'h72b6] <= 8'h1;
		memory[16'h72b7] <= 8'hb3;
		memory[16'h72b8] <= 8'hba;
		memory[16'h72b9] <= 8'he3;
		memory[16'h72ba] <= 8'h3d;
		memory[16'h72bb] <= 8'h98;
		memory[16'h72bc] <= 8'h9b;
		memory[16'h72bd] <= 8'h4e;
		memory[16'h72be] <= 8'h84;
		memory[16'h72bf] <= 8'h1b;
		memory[16'h72c0] <= 8'h55;
		memory[16'h72c1] <= 8'hfb;
		memory[16'h72c2] <= 8'h54;
		memory[16'h72c3] <= 8'hca;
		memory[16'h72c4] <= 8'hdb;
		memory[16'h72c5] <= 8'hdc;
		memory[16'h72c6] <= 8'h21;
		memory[16'h72c7] <= 8'h4b;
		memory[16'h72c8] <= 8'he4;
		memory[16'h72c9] <= 8'h68;
		memory[16'h72ca] <= 8'h5c;
		memory[16'h72cb] <= 8'hbe;
		memory[16'h72cc] <= 8'h6c;
		memory[16'h72cd] <= 8'ha8;
		memory[16'h72ce] <= 8'hbd;
		memory[16'h72cf] <= 8'h2a;
		memory[16'h72d0] <= 8'h2c;
		memory[16'h72d1] <= 8'h60;
		memory[16'h72d2] <= 8'h53;
		memory[16'h72d3] <= 8'hec;
		memory[16'h72d4] <= 8'h76;
		memory[16'h72d5] <= 8'h54;
		memory[16'h72d6] <= 8'h9f;
		memory[16'h72d7] <= 8'h30;
		memory[16'h72d8] <= 8'h37;
		memory[16'h72d9] <= 8'hdc;
		memory[16'h72da] <= 8'hc8;
		memory[16'h72db] <= 8'hd3;
		memory[16'h72dc] <= 8'h2b;
		memory[16'h72dd] <= 8'h4d;
		memory[16'h72de] <= 8'hee;
		memory[16'h72df] <= 8'h80;
		memory[16'h72e0] <= 8'h48;
		memory[16'h72e1] <= 8'h43;
		memory[16'h72e2] <= 8'h4a;
		memory[16'h72e3] <= 8'h23;
		memory[16'h72e4] <= 8'h1f;
		memory[16'h72e5] <= 8'h6b;
		memory[16'h72e6] <= 8'h6e;
		memory[16'h72e7] <= 8'h3;
		memory[16'h72e8] <= 8'hd3;
		memory[16'h72e9] <= 8'hca;
		memory[16'h72ea] <= 8'hc2;
		memory[16'h72eb] <= 8'h3f;
		memory[16'h72ec] <= 8'h72;
		memory[16'h72ed] <= 8'h7f;
		memory[16'h72ee] <= 8'h6a;
		memory[16'h72ef] <= 8'h9e;
		memory[16'h72f0] <= 8'hdf;
		memory[16'h72f1] <= 8'hbd;
		memory[16'h72f2] <= 8'h8a;
		memory[16'h72f3] <= 8'h55;
		memory[16'h72f4] <= 8'h12;
		memory[16'h72f5] <= 8'h29;
		memory[16'h72f6] <= 8'h85;
		memory[16'h72f7] <= 8'h49;
		memory[16'h72f8] <= 8'h6;
		memory[16'h72f9] <= 8'h4e;
		memory[16'h72fa] <= 8'h1c;
		memory[16'h72fb] <= 8'h31;
		memory[16'h72fc] <= 8'h9b;
		memory[16'h72fd] <= 8'hb;
		memory[16'h72fe] <= 8'hb1;
		memory[16'h72ff] <= 8'he3;
		memory[16'h7300] <= 8'h4e;
		memory[16'h7301] <= 8'hfb;
		memory[16'h7302] <= 8'h7;
		memory[16'h7303] <= 8'h6d;
		memory[16'h7304] <= 8'h67;
		memory[16'h7305] <= 8'h75;
		memory[16'h7306] <= 8'h71;
		memory[16'h7307] <= 8'h3a;
		memory[16'h7308] <= 8'h40;
		memory[16'h7309] <= 8'h33;
		memory[16'h730a] <= 8'h7a;
		memory[16'h730b] <= 8'hb2;
		memory[16'h730c] <= 8'hb2;
		memory[16'h730d] <= 8'he4;
		memory[16'h730e] <= 8'h51;
		memory[16'h730f] <= 8'h92;
		memory[16'h7310] <= 8'ha1;
		memory[16'h7311] <= 8'hdb;
		memory[16'h7312] <= 8'he7;
		memory[16'h7313] <= 8'hb3;
		memory[16'h7314] <= 8'h5;
		memory[16'h7315] <= 8'h6d;
		memory[16'h7316] <= 8'hfd;
		memory[16'h7317] <= 8'hb;
		memory[16'h7318] <= 8'hbb;
		memory[16'h7319] <= 8'h19;
		memory[16'h731a] <= 8'h3c;
		memory[16'h731b] <= 8'h56;
		memory[16'h731c] <= 8'h24;
		memory[16'h731d] <= 8'hed;
		memory[16'h731e] <= 8'h39;
		memory[16'h731f] <= 8'h72;
		memory[16'h7320] <= 8'he8;
		memory[16'h7321] <= 8'h40;
		memory[16'h7322] <= 8'he0;
		memory[16'h7323] <= 8'h4f;
		memory[16'h7324] <= 8'hb6;
		memory[16'h7325] <= 8'h51;
		memory[16'h7326] <= 8'h8a;
		memory[16'h7327] <= 8'hf6;
		memory[16'h7328] <= 8'h84;
		memory[16'h7329] <= 8'h4;
		memory[16'h732a] <= 8'ha8;
		memory[16'h732b] <= 8'h36;
		memory[16'h732c] <= 8'he8;
		memory[16'h732d] <= 8'hf9;
		memory[16'h732e] <= 8'hc8;
		memory[16'h732f] <= 8'h89;
		memory[16'h7330] <= 8'hd5;
		memory[16'h7331] <= 8'hb0;
		memory[16'h7332] <= 8'h3d;
		memory[16'h7333] <= 8'hda;
		memory[16'h7334] <= 8'h1d;
		memory[16'h7335] <= 8'h3a;
		memory[16'h7336] <= 8'he5;
		memory[16'h7337] <= 8'hd8;
		memory[16'h7338] <= 8'h53;
		memory[16'h7339] <= 8'h21;
		memory[16'h733a] <= 8'h2e;
		memory[16'h733b] <= 8'h78;
		memory[16'h733c] <= 8'he;
		memory[16'h733d] <= 8'h67;
		memory[16'h733e] <= 8'hea;
		memory[16'h733f] <= 8'hf6;
		memory[16'h7340] <= 8'ha8;
		memory[16'h7341] <= 8'hca;
		memory[16'h7342] <= 8'h46;
		memory[16'h7343] <= 8'h5e;
		memory[16'h7344] <= 8'h1b;
		memory[16'h7345] <= 8'hd0;
		memory[16'h7346] <= 8'h54;
		memory[16'h7347] <= 8'h9f;
		memory[16'h7348] <= 8'hd4;
		memory[16'h7349] <= 8'hfc;
		memory[16'h734a] <= 8'hd6;
		memory[16'h734b] <= 8'hbc;
		memory[16'h734c] <= 8'hf6;
		memory[16'h734d] <= 8'h9e;
		memory[16'h734e] <= 8'h45;
		memory[16'h734f] <= 8'hcb;
		memory[16'h7350] <= 8'h4e;
		memory[16'h7351] <= 8'h82;
		memory[16'h7352] <= 8'ha5;
		memory[16'h7353] <= 8'h6b;
		memory[16'h7354] <= 8'hbc;
		memory[16'h7355] <= 8'h8a;
		memory[16'h7356] <= 8'h43;
		memory[16'h7357] <= 8'h10;
		memory[16'h7358] <= 8'hab;
		memory[16'h7359] <= 8'h71;
		memory[16'h735a] <= 8'h88;
		memory[16'h735b] <= 8'hb9;
		memory[16'h735c] <= 8'hd9;
		memory[16'h735d] <= 8'h72;
		memory[16'h735e] <= 8'haf;
		memory[16'h735f] <= 8'h81;
		memory[16'h7360] <= 8'h3d;
		memory[16'h7361] <= 8'hf5;
		memory[16'h7362] <= 8'hdf;
		memory[16'h7363] <= 8'h58;
		memory[16'h7364] <= 8'hc5;
		memory[16'h7365] <= 8'h33;
		memory[16'h7366] <= 8'hf8;
		memory[16'h7367] <= 8'h99;
		memory[16'h7368] <= 8'h2f;
		memory[16'h7369] <= 8'hce;
		memory[16'h736a] <= 8'h55;
		memory[16'h736b] <= 8'h25;
		memory[16'h736c] <= 8'h6c;
		memory[16'h736d] <= 8'h9b;
		memory[16'h736e] <= 8'hf0;
		memory[16'h736f] <= 8'hbb;
		memory[16'h7370] <= 8'h1d;
		memory[16'h7371] <= 8'h95;
		memory[16'h7372] <= 8'h26;
		memory[16'h7373] <= 8'hda;
		memory[16'h7374] <= 8'h1f;
		memory[16'h7375] <= 8'h6a;
		memory[16'h7376] <= 8'hea;
		memory[16'h7377] <= 8'hca;
		memory[16'h7378] <= 8'hdb;
		memory[16'h7379] <= 8'h72;
		memory[16'h737a] <= 8'h83;
		memory[16'h737b] <= 8'hb4;
		memory[16'h737c] <= 8'he4;
		memory[16'h737d] <= 8'h33;
		memory[16'h737e] <= 8'h35;
		memory[16'h737f] <= 8'h21;
		memory[16'h7380] <= 8'h28;
		memory[16'h7381] <= 8'h14;
		memory[16'h7382] <= 8'h7a;
		memory[16'h7383] <= 8'hee;
		memory[16'h7384] <= 8'h47;
		memory[16'h7385] <= 8'h72;
		memory[16'h7386] <= 8'h87;
		memory[16'h7387] <= 8'h77;
		memory[16'h7388] <= 8'h40;
		memory[16'h7389] <= 8'hdd;
		memory[16'h738a] <= 8'h9c;
		memory[16'h738b] <= 8'hac;
		memory[16'h738c] <= 8'h78;
		memory[16'h738d] <= 8'h8d;
		memory[16'h738e] <= 8'h67;
		memory[16'h738f] <= 8'h95;
		memory[16'h7390] <= 8'h22;
		memory[16'h7391] <= 8'h8e;
		memory[16'h7392] <= 8'h6f;
		memory[16'h7393] <= 8'h42;
		memory[16'h7394] <= 8'hf8;
		memory[16'h7395] <= 8'h59;
		memory[16'h7396] <= 8'hc;
		memory[16'h7397] <= 8'hd3;
		memory[16'h7398] <= 8'hcb;
		memory[16'h7399] <= 8'h90;
		memory[16'h739a] <= 8'h88;
		memory[16'h739b] <= 8'hb0;
		memory[16'h739c] <= 8'hc3;
		memory[16'h739d] <= 8'hbd;
		memory[16'h739e] <= 8'hd1;
		memory[16'h739f] <= 8'heb;
		memory[16'h73a0] <= 8'hd2;
		memory[16'h73a1] <= 8'h4b;
		memory[16'h73a2] <= 8'hd9;
		memory[16'h73a3] <= 8'h19;
		memory[16'h73a4] <= 8'hbd;
		memory[16'h73a5] <= 8'h61;
		memory[16'h73a6] <= 8'h90;
		memory[16'h73a7] <= 8'hfd;
		memory[16'h73a8] <= 8'h3e;
		memory[16'h73a9] <= 8'h2d;
		memory[16'h73aa] <= 8'haa;
		memory[16'h73ab] <= 8'hb6;
		memory[16'h73ac] <= 8'hba;
		memory[16'h73ad] <= 8'h11;
		memory[16'h73ae] <= 8'h4b;
		memory[16'h73af] <= 8'hdc;
		memory[16'h73b0] <= 8'h9f;
		memory[16'h73b1] <= 8'hbb;
		memory[16'h73b2] <= 8'h1e;
		memory[16'h73b3] <= 8'h97;
		memory[16'h73b4] <= 8'h14;
		memory[16'h73b5] <= 8'h2b;
		memory[16'h73b6] <= 8'h6b;
		memory[16'h73b7] <= 8'he0;
		memory[16'h73b8] <= 8'hbb;
		memory[16'h73b9] <= 8'hf3;
		memory[16'h73ba] <= 8'h90;
		memory[16'h73bb] <= 8'h7e;
		memory[16'h73bc] <= 8'hb0;
		memory[16'h73bd] <= 8'h61;
		memory[16'h73be] <= 8'h69;
		memory[16'h73bf] <= 8'h82;
		memory[16'h73c0] <= 8'had;
		memory[16'h73c1] <= 8'h43;
		memory[16'h73c2] <= 8'h9c;
		memory[16'h73c3] <= 8'h6a;
		memory[16'h73c4] <= 8'ha4;
		memory[16'h73c5] <= 8'h2c;
		memory[16'h73c6] <= 8'h68;
		memory[16'h73c7] <= 8'he2;
		memory[16'h73c8] <= 8'h59;
		memory[16'h73c9] <= 8'h12;
		memory[16'h73ca] <= 8'h98;
		memory[16'h73cb] <= 8'h13;
		memory[16'h73cc] <= 8'h23;
		memory[16'h73cd] <= 8'he3;
		memory[16'h73ce] <= 8'hf0;
		memory[16'h73cf] <= 8'hc3;
		memory[16'h73d0] <= 8'h9e;
		memory[16'h73d1] <= 8'he;
		memory[16'h73d2] <= 8'h5a;
		memory[16'h73d3] <= 8'hb3;
		memory[16'h73d4] <= 8'h39;
		memory[16'h73d5] <= 8'hc5;
		memory[16'h73d6] <= 8'h93;
		memory[16'h73d7] <= 8'hf4;
		memory[16'h73d8] <= 8'hb8;
		memory[16'h73d9] <= 8'h23;
		memory[16'h73da] <= 8'h72;
		memory[16'h73db] <= 8'h69;
		memory[16'h73dc] <= 8'h84;
		memory[16'h73dd] <= 8'hdc;
		memory[16'h73de] <= 8'heb;
		memory[16'h73df] <= 8'h31;
		memory[16'h73e0] <= 8'h1f;
		memory[16'h73e1] <= 8'h87;
		memory[16'h73e2] <= 8'h9c;
		memory[16'h73e3] <= 8'hc3;
		memory[16'h73e4] <= 8'hb4;
		memory[16'h73e5] <= 8'h4;
		memory[16'h73e6] <= 8'ha5;
		memory[16'h73e7] <= 8'hd;
		memory[16'h73e8] <= 8'h16;
		memory[16'h73e9] <= 8'h3d;
		memory[16'h73ea] <= 8'h21;
		memory[16'h73eb] <= 8'h39;
		memory[16'h73ec] <= 8'h20;
		memory[16'h73ed] <= 8'h11;
		memory[16'h73ee] <= 8'hfc;
		memory[16'h73ef] <= 8'hbf;
		memory[16'h73f0] <= 8'h1f;
		memory[16'h73f1] <= 8'h57;
		memory[16'h73f2] <= 8'h72;
		memory[16'h73f3] <= 8'h59;
		memory[16'h73f4] <= 8'h1c;
		memory[16'h73f5] <= 8'h5;
		memory[16'h73f6] <= 8'h4d;
		memory[16'h73f7] <= 8'hd5;
		memory[16'h73f8] <= 8'h28;
		memory[16'h73f9] <= 8'hc0;
		memory[16'h73fa] <= 8'h3e;
		memory[16'h73fb] <= 8'hac;
		memory[16'h73fc] <= 8'h9c;
		memory[16'h73fd] <= 8'h29;
		memory[16'h73fe] <= 8'hde;
		memory[16'h73ff] <= 8'hbb;
		memory[16'h7400] <= 8'hb1;
		memory[16'h7401] <= 8'h7a;
		memory[16'h7402] <= 8'h7e;
		memory[16'h7403] <= 8'h65;
		memory[16'h7404] <= 8'h7e;
		memory[16'h7405] <= 8'h23;
		memory[16'h7406] <= 8'h72;
		memory[16'h7407] <= 8'h94;
		memory[16'h7408] <= 8'h60;
		memory[16'h7409] <= 8'h93;
		memory[16'h740a] <= 8'hcd;
		memory[16'h740b] <= 8'h80;
		memory[16'h740c] <= 8'ha4;
		memory[16'h740d] <= 8'hca;
		memory[16'h740e] <= 8'h3f;
		memory[16'h740f] <= 8'hc4;
		memory[16'h7410] <= 8'h21;
		memory[16'h7411] <= 8'hb1;
		memory[16'h7412] <= 8'h1d;
		memory[16'h7413] <= 8'h3d;
		memory[16'h7414] <= 8'hb6;
		memory[16'h7415] <= 8'h6a;
		memory[16'h7416] <= 8'h12;
		memory[16'h7417] <= 8'hde;
		memory[16'h7418] <= 8'h2a;
		memory[16'h7419] <= 8'h50;
		memory[16'h741a] <= 8'h8b;
		memory[16'h741b] <= 8'hc6;
		memory[16'h741c] <= 8'h7a;
		memory[16'h741d] <= 8'h69;
		memory[16'h741e] <= 8'h81;
		memory[16'h741f] <= 8'h2b;
		memory[16'h7420] <= 8'he3;
		memory[16'h7421] <= 8'hff;
		memory[16'h7422] <= 8'h90;
		memory[16'h7423] <= 8'h61;
		memory[16'h7424] <= 8'h22;
		memory[16'h7425] <= 8'h2;
		memory[16'h7426] <= 8'hf5;
		memory[16'h7427] <= 8'h82;
		memory[16'h7428] <= 8'h96;
		memory[16'h7429] <= 8'hc2;
		memory[16'h742a] <= 8'h3;
		memory[16'h742b] <= 8'h3a;
		memory[16'h742c] <= 8'h8c;
		memory[16'h742d] <= 8'h42;
		memory[16'h742e] <= 8'hfe;
		memory[16'h742f] <= 8'had;
		memory[16'h7430] <= 8'hf4;
		memory[16'h7431] <= 8'h1b;
		memory[16'h7432] <= 8'heb;
		memory[16'h7433] <= 8'haa;
		memory[16'h7434] <= 8'h86;
		memory[16'h7435] <= 8'hfd;
		memory[16'h7436] <= 8'h89;
		memory[16'h7437] <= 8'hb0;
		memory[16'h7438] <= 8'h4e;
		memory[16'h7439] <= 8'h14;
		memory[16'h743a] <= 8'h77;
		memory[16'h743b] <= 8'hc8;
		memory[16'h743c] <= 8'h7d;
		memory[16'h743d] <= 8'hf8;
		memory[16'h743e] <= 8'hf3;
		memory[16'h743f] <= 8'h60;
		memory[16'h7440] <= 8'hf8;
		memory[16'h7441] <= 8'h83;
		memory[16'h7442] <= 8'hc1;
		memory[16'h7443] <= 8'h1a;
		memory[16'h7444] <= 8'h85;
		memory[16'h7445] <= 8'hb6;
		memory[16'h7446] <= 8'h9d;
		memory[16'h7447] <= 8'h1b;
		memory[16'h7448] <= 8'h78;
		memory[16'h7449] <= 8'ha0;
		memory[16'h744a] <= 8'h56;
		memory[16'h744b] <= 8'h5;
		memory[16'h744c] <= 8'he2;
		memory[16'h744d] <= 8'h54;
		memory[16'h744e] <= 8'hb2;
		memory[16'h744f] <= 8'hd6;
		memory[16'h7450] <= 8'h70;
		memory[16'h7451] <= 8'h9d;
		memory[16'h7452] <= 8'h81;
		memory[16'h7453] <= 8'hf6;
		memory[16'h7454] <= 8'h9b;
		memory[16'h7455] <= 8'ha;
		memory[16'h7456] <= 8'ha6;
		memory[16'h7457] <= 8'he9;
		memory[16'h7458] <= 8'h1e;
		memory[16'h7459] <= 8'h1d;
		memory[16'h745a] <= 8'hb1;
		memory[16'h745b] <= 8'h9b;
		memory[16'h745c] <= 8'h16;
		memory[16'h745d] <= 8'ha4;
		memory[16'h745e] <= 8'hfb;
		memory[16'h745f] <= 8'he;
		memory[16'h7460] <= 8'h27;
		memory[16'h7461] <= 8'hbc;
		memory[16'h7462] <= 8'h28;
		memory[16'h7463] <= 8'hac;
		memory[16'h7464] <= 8'h72;
		memory[16'h7465] <= 8'hc5;
		memory[16'h7466] <= 8'hc8;
		memory[16'h7467] <= 8'hea;
		memory[16'h7468] <= 8'h65;
		memory[16'h7469] <= 8'h1e;
		memory[16'h746a] <= 8'hef;
		memory[16'h746b] <= 8'h48;
		memory[16'h746c] <= 8'h72;
		memory[16'h746d] <= 8'ha2;
		memory[16'h746e] <= 8'h1e;
		memory[16'h746f] <= 8'he2;
		memory[16'h7470] <= 8'h3f;
		memory[16'h7471] <= 8'h9f;
		memory[16'h7472] <= 8'hd8;
		memory[16'h7473] <= 8'hda;
		memory[16'h7474] <= 8'ha9;
		memory[16'h7475] <= 8'h7f;
		memory[16'h7476] <= 8'hc3;
		memory[16'h7477] <= 8'hc7;
		memory[16'h7478] <= 8'h9c;
		memory[16'h7479] <= 8'h74;
		memory[16'h747a] <= 8'h62;
		memory[16'h747b] <= 8'hb2;
		memory[16'h747c] <= 8'h18;
		memory[16'h747d] <= 8'h5d;
		memory[16'h747e] <= 8'hc0;
		memory[16'h747f] <= 8'h3f;
		memory[16'h7480] <= 8'h19;
		memory[16'h7481] <= 8'he9;
		memory[16'h7482] <= 8'hec;
		memory[16'h7483] <= 8'h8b;
		memory[16'h7484] <= 8'hae;
		memory[16'h7485] <= 8'hb4;
		memory[16'h7486] <= 8'h76;
		memory[16'h7487] <= 8'h14;
		memory[16'h7488] <= 8'hd2;
		memory[16'h7489] <= 8'h65;
		memory[16'h748a] <= 8'h5c;
		memory[16'h748b] <= 8'h44;
		memory[16'h748c] <= 8'h7;
		memory[16'h748d] <= 8'h7a;
		memory[16'h748e] <= 8'h27;
		memory[16'h748f] <= 8'h47;
		memory[16'h7490] <= 8'h1a;
		memory[16'h7491] <= 8'hff;
		memory[16'h7492] <= 8'h21;
		memory[16'h7493] <= 8'hc3;
		memory[16'h7494] <= 8'h7e;
		memory[16'h7495] <= 8'he5;
		memory[16'h7496] <= 8'h8b;
		memory[16'h7497] <= 8'h1b;
		memory[16'h7498] <= 8'h59;
		memory[16'h7499] <= 8'hed;
		memory[16'h749a] <= 8'hcd;
		memory[16'h749b] <= 8'h72;
		memory[16'h749c] <= 8'h4b;
		memory[16'h749d] <= 8'h8e;
		memory[16'h749e] <= 8'hb1;
		memory[16'h749f] <= 8'h64;
		memory[16'h74a0] <= 8'h77;
		memory[16'h74a1] <= 8'h9d;
		memory[16'h74a2] <= 8'hf0;
		memory[16'h74a3] <= 8'h25;
		memory[16'h74a4] <= 8'h51;
		memory[16'h74a5] <= 8'h66;
		memory[16'h74a6] <= 8'h39;
		memory[16'h74a7] <= 8'h23;
		memory[16'h74a8] <= 8'hcb;
		memory[16'h74a9] <= 8'h95;
		memory[16'h74aa] <= 8'h68;
		memory[16'h74ab] <= 8'hd3;
		memory[16'h74ac] <= 8'h10;
		memory[16'h74ad] <= 8'h8f;
		memory[16'h74ae] <= 8'h1a;
		memory[16'h74af] <= 8'h2a;
		memory[16'h74b0] <= 8'h8e;
		memory[16'h74b1] <= 8'h3b;
		memory[16'h74b2] <= 8'hed;
		memory[16'h74b3] <= 8'hd;
		memory[16'h74b4] <= 8'h20;
		memory[16'h74b5] <= 8'h78;
		memory[16'h74b6] <= 8'h28;
		memory[16'h74b7] <= 8'h7a;
		memory[16'h74b8] <= 8'h66;
		memory[16'h74b9] <= 8'hf5;
		memory[16'h74ba] <= 8'hec;
		memory[16'h74bb] <= 8'hb1;
		memory[16'h74bc] <= 8'h83;
		memory[16'h74bd] <= 8'h9d;
		memory[16'h74be] <= 8'h15;
		memory[16'h74bf] <= 8'hfa;
		memory[16'h74c0] <= 8'h3b;
		memory[16'h74c1] <= 8'h5;
		memory[16'h74c2] <= 8'h20;
		memory[16'h74c3] <= 8'h8c;
		memory[16'h74c4] <= 8'h6b;
		memory[16'h74c5] <= 8'h59;
		memory[16'h74c6] <= 8'hb0;
		memory[16'h74c7] <= 8'h37;
		memory[16'h74c8] <= 8'hef;
		memory[16'h74c9] <= 8'h18;
		memory[16'h74ca] <= 8'ha;
		memory[16'h74cb] <= 8'hff;
		memory[16'h74cc] <= 8'ha7;
		memory[16'h74cd] <= 8'h24;
		memory[16'h74ce] <= 8'h29;
		memory[16'h74cf] <= 8'h35;
		memory[16'h74d0] <= 8'h5f;
		memory[16'h74d1] <= 8'h16;
		memory[16'h74d2] <= 8'h42;
		memory[16'h74d3] <= 8'h80;
		memory[16'h74d4] <= 8'h8f;
		memory[16'h74d5] <= 8'h6a;
		memory[16'h74d6] <= 8'hfa;
		memory[16'h74d7] <= 8'hf5;
		memory[16'h74d8] <= 8'h60;
		memory[16'h74d9] <= 8'he6;
		memory[16'h74da] <= 8'ha6;
		memory[16'h74db] <= 8'he3;
		memory[16'h74dc] <= 8'h83;
		memory[16'h74dd] <= 8'hbb;
		memory[16'h74de] <= 8'hde;
		memory[16'h74df] <= 8'hbe;
		memory[16'h74e0] <= 8'hc1;
		memory[16'h74e1] <= 8'hfe;
		memory[16'h74e2] <= 8'h4b;
		memory[16'h74e3] <= 8'h2c;
		memory[16'h74e4] <= 8'h57;
		memory[16'h74e5] <= 8'hfb;
		memory[16'h74e6] <= 8'h63;
		memory[16'h74e7] <= 8'h46;
		memory[16'h74e8] <= 8'h13;
		memory[16'h74e9] <= 8'h6d;
		memory[16'h74ea] <= 8'h45;
		memory[16'h74eb] <= 8'hba;
		memory[16'h74ec] <= 8'h91;
		memory[16'h74ed] <= 8'h6e;
		memory[16'h74ee] <= 8'hef;
		memory[16'h74ef] <= 8'hf1;
		memory[16'h74f0] <= 8'h85;
		memory[16'h74f1] <= 8'h32;
		memory[16'h74f2] <= 8'h71;
		memory[16'h74f3] <= 8'h14;
		memory[16'h74f4] <= 8'h9c;
		memory[16'h74f5] <= 8'h6b;
		memory[16'h74f6] <= 8'h9;
		memory[16'h74f7] <= 8'hfc;
		memory[16'h74f8] <= 8'h51;
		memory[16'h74f9] <= 8'haf;
		memory[16'h74fa] <= 8'he0;
		memory[16'h74fb] <= 8'hd4;
		memory[16'h74fc] <= 8'h6a;
		memory[16'h74fd] <= 8'hbe;
		memory[16'h74fe] <= 8'h93;
		memory[16'h74ff] <= 8'h2b;
		memory[16'h7500] <= 8'hbc;
		memory[16'h7501] <= 8'hde;
		memory[16'h7502] <= 8'h58;
		memory[16'h7503] <= 8'h13;
		memory[16'h7504] <= 8'hd9;
		memory[16'h7505] <= 8'hbb;
		memory[16'h7506] <= 8'h5a;
		memory[16'h7507] <= 8'hec;
		memory[16'h7508] <= 8'h29;
		memory[16'h7509] <= 8'h9f;
		memory[16'h750a] <= 8'ha6;
		memory[16'h750b] <= 8'hba;
		memory[16'h750c] <= 8'he;
		memory[16'h750d] <= 8'h95;
		memory[16'h750e] <= 8'hab;
		memory[16'h750f] <= 8'h93;
		memory[16'h7510] <= 8'hc7;
		memory[16'h7511] <= 8'h1c;
		memory[16'h7512] <= 8'ha7;
		memory[16'h7513] <= 8'h64;
		memory[16'h7514] <= 8'h87;
		memory[16'h7515] <= 8'hb0;
		memory[16'h7516] <= 8'h60;
		memory[16'h7517] <= 8'hd8;
		memory[16'h7518] <= 8'h5f;
		memory[16'h7519] <= 8'h40;
		memory[16'h751a] <= 8'had;
		memory[16'h751b] <= 8'hc9;
		memory[16'h751c] <= 8'hfe;
		memory[16'h751d] <= 8'h40;
		memory[16'h751e] <= 8'hf5;
		memory[16'h751f] <= 8'hba;
		memory[16'h7520] <= 8'h1e;
		memory[16'h7521] <= 8'h4d;
		memory[16'h7522] <= 8'hce;
		memory[16'h7523] <= 8'hf7;
		memory[16'h7524] <= 8'h8;
		memory[16'h7525] <= 8'h28;
		memory[16'h7526] <= 8'he3;
		memory[16'h7527] <= 8'h31;
		memory[16'h7528] <= 8'hc7;
		memory[16'h7529] <= 8'h89;
		memory[16'h752a] <= 8'hec;
		memory[16'h752b] <= 8'hd5;
		memory[16'h752c] <= 8'h1e;
		memory[16'h752d] <= 8'h97;
		memory[16'h752e] <= 8'h68;
		memory[16'h752f] <= 8'he6;
		memory[16'h7530] <= 8'hb4;
		memory[16'h7531] <= 8'hf;
		memory[16'h7532] <= 8'h4a;
		memory[16'h7533] <= 8'h3b;
		memory[16'h7534] <= 8'hbf;
		memory[16'h7535] <= 8'haa;
		memory[16'h7536] <= 8'h14;
		memory[16'h7537] <= 8'h1e;
		memory[16'h7538] <= 8'heb;
		memory[16'h7539] <= 8'hc1;
		memory[16'h753a] <= 8'he8;
		memory[16'h753b] <= 8'he9;
		memory[16'h753c] <= 8'h1;
		memory[16'h753d] <= 8'hdd;
		memory[16'h753e] <= 8'ha4;
		memory[16'h753f] <= 8'h1f;
		memory[16'h7540] <= 8'h2a;
		memory[16'h7541] <= 8'h72;
		memory[16'h7542] <= 8'h16;
		memory[16'h7543] <= 8'h32;
		memory[16'h7544] <= 8'h9a;
		memory[16'h7545] <= 8'hf9;
		memory[16'h7546] <= 8'h64;
		memory[16'h7547] <= 8'h61;
		memory[16'h7548] <= 8'h82;
		memory[16'h7549] <= 8'h50;
		memory[16'h754a] <= 8'h37;
		memory[16'h754b] <= 8'ha0;
		memory[16'h754c] <= 8'he7;
		memory[16'h754d] <= 8'h9f;
		memory[16'h754e] <= 8'h86;
		memory[16'h754f] <= 8'h9b;
		memory[16'h7550] <= 8'haf;
		memory[16'h7551] <= 8'hd0;
		memory[16'h7552] <= 8'hd7;
		memory[16'h7553] <= 8'h6e;
		memory[16'h7554] <= 8'h7b;
		memory[16'h7555] <= 8'heb;
		memory[16'h7556] <= 8'h8d;
		memory[16'h7557] <= 8'h66;
		memory[16'h7558] <= 8'hac;
		memory[16'h7559] <= 8'h75;
		memory[16'h755a] <= 8'h4f;
		memory[16'h755b] <= 8'had;
		memory[16'h755c] <= 8'h52;
		memory[16'h755d] <= 8'hf3;
		memory[16'h755e] <= 8'hcc;
		memory[16'h755f] <= 8'h7c;
		memory[16'h7560] <= 8'h65;
		memory[16'h7561] <= 8'he2;
		memory[16'h7562] <= 8'hae;
		memory[16'h7563] <= 8'hff;
		memory[16'h7564] <= 8'hdb;
		memory[16'h7565] <= 8'h12;
		memory[16'h7566] <= 8'h61;
		memory[16'h7567] <= 8'h5d;
		memory[16'h7568] <= 8'h62;
		memory[16'h7569] <= 8'h98;
		memory[16'h756a] <= 8'hfd;
		memory[16'h756b] <= 8'h4a;
		memory[16'h756c] <= 8'h37;
		memory[16'h756d] <= 8'h84;
		memory[16'h756e] <= 8'he5;
		memory[16'h756f] <= 8'he6;
		memory[16'h7570] <= 8'h54;
		memory[16'h7571] <= 8'hbc;
		memory[16'h7572] <= 8'h55;
		memory[16'h7573] <= 8'hcf;
		memory[16'h7574] <= 8'ha7;
		memory[16'h7575] <= 8'he2;
		memory[16'h7576] <= 8'h35;
		memory[16'h7577] <= 8'h53;
		memory[16'h7578] <= 8'h57;
		memory[16'h7579] <= 8'h85;
		memory[16'h757a] <= 8'h0;
		memory[16'h757b] <= 8'ha9;
		memory[16'h757c] <= 8'h78;
		memory[16'h757d] <= 8'hcc;
		memory[16'h757e] <= 8'h25;
		memory[16'h757f] <= 8'hde;
		memory[16'h7580] <= 8'hae;
		memory[16'h7581] <= 8'hd3;
		memory[16'h7582] <= 8'hdd;
		memory[16'h7583] <= 8'h89;
		memory[16'h7584] <= 8'he6;
		memory[16'h7585] <= 8'h3e;
		memory[16'h7586] <= 8'he6;
		memory[16'h7587] <= 8'h48;
		memory[16'h7588] <= 8'hd6;
		memory[16'h7589] <= 8'he4;
		memory[16'h758a] <= 8'h92;
		memory[16'h758b] <= 8'he;
		memory[16'h758c] <= 8'h68;
		memory[16'h758d] <= 8'h78;
		memory[16'h758e] <= 8'hf4;
		memory[16'h758f] <= 8'hbc;
		memory[16'h7590] <= 8'h34;
		memory[16'h7591] <= 8'h49;
		memory[16'h7592] <= 8'h8c;
		memory[16'h7593] <= 8'hdc;
		memory[16'h7594] <= 8'h2b;
		memory[16'h7595] <= 8'hc1;
		memory[16'h7596] <= 8'h2f;
		memory[16'h7597] <= 8'h82;
		memory[16'h7598] <= 8'h46;
		memory[16'h7599] <= 8'h30;
		memory[16'h759a] <= 8'h2b;
		memory[16'h759b] <= 8'hbf;
		memory[16'h759c] <= 8'hfc;
		memory[16'h759d] <= 8'h50;
		memory[16'h759e] <= 8'h9d;
		memory[16'h759f] <= 8'hab;
		memory[16'h75a0] <= 8'h24;
		memory[16'h75a1] <= 8'h7a;
		memory[16'h75a2] <= 8'h34;
		memory[16'h75a3] <= 8'ha;
		memory[16'h75a4] <= 8'hb9;
		memory[16'h75a5] <= 8'h1b;
		memory[16'h75a6] <= 8'h52;
		memory[16'h75a7] <= 8'h8f;
		memory[16'h75a8] <= 8'hff;
		memory[16'h75a9] <= 8'he5;
		memory[16'h75aa] <= 8'h9d;
		memory[16'h75ab] <= 8'h67;
		memory[16'h75ac] <= 8'h5d;
		memory[16'h75ad] <= 8'h92;
		memory[16'h75ae] <= 8'h23;
		memory[16'h75af] <= 8'h91;
		memory[16'h75b0] <= 8'hdb;
		memory[16'h75b1] <= 8'haf;
		memory[16'h75b2] <= 8'h6d;
		memory[16'h75b3] <= 8'h7;
		memory[16'h75b4] <= 8'h71;
		memory[16'h75b5] <= 8'h9d;
		memory[16'h75b6] <= 8'h89;
		memory[16'h75b7] <= 8'hb7;
		memory[16'h75b8] <= 8'hcd;
		memory[16'h75b9] <= 8'hb5;
		memory[16'h75ba] <= 8'h76;
		memory[16'h75bb] <= 8'hc9;
		memory[16'h75bc] <= 8'h5;
		memory[16'h75bd] <= 8'h13;
		memory[16'h75be] <= 8'h74;
		memory[16'h75bf] <= 8'h29;
		memory[16'h75c0] <= 8'h8e;
		memory[16'h75c1] <= 8'ha9;
		memory[16'h75c2] <= 8'h33;
		memory[16'h75c3] <= 8'h47;
		memory[16'h75c4] <= 8'hc4;
		memory[16'h75c5] <= 8'h86;
		memory[16'h75c6] <= 8'hd6;
		memory[16'h75c7] <= 8'hc3;
		memory[16'h75c8] <= 8'h6b;
		memory[16'h75c9] <= 8'h74;
		memory[16'h75ca] <= 8'h2a;
		memory[16'h75cb] <= 8'hc8;
		memory[16'h75cc] <= 8'h6;
		memory[16'h75cd] <= 8'h4d;
		memory[16'h75ce] <= 8'h59;
		memory[16'h75cf] <= 8'he1;
		memory[16'h75d0] <= 8'hfd;
		memory[16'h75d1] <= 8'hc7;
		memory[16'h75d2] <= 8'he8;
		memory[16'h75d3] <= 8'h6e;
		memory[16'h75d4] <= 8'h64;
		memory[16'h75d5] <= 8'h72;
		memory[16'h75d6] <= 8'h25;
		memory[16'h75d7] <= 8'h31;
		memory[16'h75d8] <= 8'h27;
		memory[16'h75d9] <= 8'h9c;
		memory[16'h75da] <= 8'hfa;
		memory[16'h75db] <= 8'h2c;
		memory[16'h75dc] <= 8'haf;
		memory[16'h75dd] <= 8'h6f;
		memory[16'h75de] <= 8'h56;
		memory[16'h75df] <= 8'h3d;
		memory[16'h75e0] <= 8'h18;
		memory[16'h75e1] <= 8'h89;
		memory[16'h75e2] <= 8'h84;
		memory[16'h75e3] <= 8'hdc;
		memory[16'h75e4] <= 8'hf;
		memory[16'h75e5] <= 8'h5b;
		memory[16'h75e6] <= 8'h9f;
		memory[16'h75e7] <= 8'h7a;
		memory[16'h75e8] <= 8'hcf;
		memory[16'h75e9] <= 8'hc9;
		memory[16'h75ea] <= 8'h42;
		memory[16'h75eb] <= 8'hd5;
		memory[16'h75ec] <= 8'h16;
		memory[16'h75ed] <= 8'h9c;
		memory[16'h75ee] <= 8'hb6;
		memory[16'h75ef] <= 8'h13;
		memory[16'h75f0] <= 8'h63;
		memory[16'h75f1] <= 8'h9f;
		memory[16'h75f2] <= 8'h81;
		memory[16'h75f3] <= 8'hc7;
		memory[16'h75f4] <= 8'h11;
		memory[16'h75f5] <= 8'ha7;
		memory[16'h75f6] <= 8'hf8;
		memory[16'h75f7] <= 8'h38;
		memory[16'h75f8] <= 8'h43;
		memory[16'h75f9] <= 8'hf2;
		memory[16'h75fa] <= 8'h64;
		memory[16'h75fb] <= 8'hf2;
		memory[16'h75fc] <= 8'h61;
		memory[16'h75fd] <= 8'hba;
		memory[16'h75fe] <= 8'h30;
		memory[16'h75ff] <= 8'h79;
		memory[16'h7600] <= 8'h44;
		memory[16'h7601] <= 8'hb4;
		memory[16'h7602] <= 8'h55;
		memory[16'h7603] <= 8'h53;
		memory[16'h7604] <= 8'hf;
		memory[16'h7605] <= 8'hf4;
		memory[16'h7606] <= 8'hce;
		memory[16'h7607] <= 8'hde;
		memory[16'h7608] <= 8'hbd;
		memory[16'h7609] <= 8'h10;
		memory[16'h760a] <= 8'hb3;
		memory[16'h760b] <= 8'hd4;
		memory[16'h760c] <= 8'hac;
		memory[16'h760d] <= 8'h6a;
		memory[16'h760e] <= 8'he7;
		memory[16'h760f] <= 8'hf;
		memory[16'h7610] <= 8'h9;
		memory[16'h7611] <= 8'h69;
		memory[16'h7612] <= 8'hd6;
		memory[16'h7613] <= 8'h1a;
		memory[16'h7614] <= 8'h10;
		memory[16'h7615] <= 8'hce;
		memory[16'h7616] <= 8'h52;
		memory[16'h7617] <= 8'h53;
		memory[16'h7618] <= 8'hc1;
		memory[16'h7619] <= 8'hb6;
		memory[16'h761a] <= 8'h45;
		memory[16'h761b] <= 8'h22;
		memory[16'h761c] <= 8'h71;
		memory[16'h761d] <= 8'h75;
		memory[16'h761e] <= 8'h9c;
		memory[16'h761f] <= 8'hb5;
		memory[16'h7620] <= 8'h2a;
		memory[16'h7621] <= 8'hf1;
		memory[16'h7622] <= 8'h8;
		memory[16'h7623] <= 8'h39;
		memory[16'h7624] <= 8'he6;
		memory[16'h7625] <= 8'hd6;
		memory[16'h7626] <= 8'h18;
		memory[16'h7627] <= 8'ha3;
		memory[16'h7628] <= 8'he7;
		memory[16'h7629] <= 8'hcb;
		memory[16'h762a] <= 8'h77;
		memory[16'h762b] <= 8'h93;
		memory[16'h762c] <= 8'h35;
		memory[16'h762d] <= 8'h5f;
		memory[16'h762e] <= 8'ha3;
		memory[16'h762f] <= 8'h3e;
		memory[16'h7630] <= 8'hc8;
		memory[16'h7631] <= 8'h79;
		memory[16'h7632] <= 8'h58;
		memory[16'h7633] <= 8'hd8;
		memory[16'h7634] <= 8'h48;
		memory[16'h7635] <= 8'haa;
		memory[16'h7636] <= 8'h2b;
		memory[16'h7637] <= 8'h9;
		memory[16'h7638] <= 8'h61;
		memory[16'h7639] <= 8'h70;
		memory[16'h763a] <= 8'h2b;
		memory[16'h763b] <= 8'hd2;
		memory[16'h763c] <= 8'he6;
		memory[16'h763d] <= 8'hc7;
		memory[16'h763e] <= 8'h87;
		memory[16'h763f] <= 8'h10;
		memory[16'h7640] <= 8'hb9;
		memory[16'h7641] <= 8'h8f;
		memory[16'h7642] <= 8'h49;
		memory[16'h7643] <= 8'h9f;
		memory[16'h7644] <= 8'h66;
		memory[16'h7645] <= 8'h61;
		memory[16'h7646] <= 8'h42;
		memory[16'h7647] <= 8'h4d;
		memory[16'h7648] <= 8'h2d;
		memory[16'h7649] <= 8'hba;
		memory[16'h764a] <= 8'he0;
		memory[16'h764b] <= 8'h62;
		memory[16'h764c] <= 8'h19;
		memory[16'h764d] <= 8'h83;
		memory[16'h764e] <= 8'ha1;
		memory[16'h764f] <= 8'he1;
		memory[16'h7650] <= 8'hfd;
		memory[16'h7651] <= 8'hf9;
		memory[16'h7652] <= 8'hb9;
		memory[16'h7653] <= 8'h45;
		memory[16'h7654] <= 8'ha4;
		memory[16'h7655] <= 8'he4;
		memory[16'h7656] <= 8'h4e;
		memory[16'h7657] <= 8'h5;
		memory[16'h7658] <= 8'h54;
		memory[16'h7659] <= 8'h79;
		memory[16'h765a] <= 8'hd7;
		memory[16'h765b] <= 8'h3a;
		memory[16'h765c] <= 8'h41;
		memory[16'h765d] <= 8'h5e;
		memory[16'h765e] <= 8'h4a;
		memory[16'h765f] <= 8'hfa;
		memory[16'h7660] <= 8'hed;
		memory[16'h7661] <= 8'h94;
		memory[16'h7662] <= 8'h99;
		memory[16'h7663] <= 8'h53;
		memory[16'h7664] <= 8'hf5;
		memory[16'h7665] <= 8'hdb;
		memory[16'h7666] <= 8'ha0;
		memory[16'h7667] <= 8'h22;
		memory[16'h7668] <= 8'h95;
		memory[16'h7669] <= 8'h81;
		memory[16'h766a] <= 8'h85;
		memory[16'h766b] <= 8'hae;
		memory[16'h766c] <= 8'h4;
		memory[16'h766d] <= 8'h26;
		memory[16'h766e] <= 8'h8f;
		memory[16'h766f] <= 8'h1;
		memory[16'h7670] <= 8'h1f;
		memory[16'h7671] <= 8'h48;
		memory[16'h7672] <= 8'h46;
		memory[16'h7673] <= 8'hc3;
		memory[16'h7674] <= 8'h2c;
		memory[16'h7675] <= 8'h94;
		memory[16'h7676] <= 8'hc8;
		memory[16'h7677] <= 8'h81;
		memory[16'h7678] <= 8'he;
		memory[16'h7679] <= 8'h9f;
		memory[16'h767a] <= 8'hbb;
		memory[16'h767b] <= 8'h4f;
		memory[16'h767c] <= 8'hfd;
		memory[16'h767d] <= 8'h6;
		memory[16'h767e] <= 8'h49;
		memory[16'h767f] <= 8'heb;
		memory[16'h7680] <= 8'h9a;
		memory[16'h7681] <= 8'he2;
		memory[16'h7682] <= 8'h3e;
		memory[16'h7683] <= 8'h8f;
		memory[16'h7684] <= 8'hbd;
		memory[16'h7685] <= 8'hdf;
		memory[16'h7686] <= 8'hb2;
		memory[16'h7687] <= 8'h53;
		memory[16'h7688] <= 8'h60;
		memory[16'h7689] <= 8'h37;
		memory[16'h768a] <= 8'h1;
		memory[16'h768b] <= 8'h64;
		memory[16'h768c] <= 8'h5d;
		memory[16'h768d] <= 8'h91;
		memory[16'h768e] <= 8'h66;
		memory[16'h768f] <= 8'h7c;
		memory[16'h7690] <= 8'hd9;
		memory[16'h7691] <= 8'hac;
		memory[16'h7692] <= 8'h40;
		memory[16'h7693] <= 8'h6;
		memory[16'h7694] <= 8'h41;
		memory[16'h7695] <= 8'h8;
		memory[16'h7696] <= 8'h87;
		memory[16'h7697] <= 8'h4f;
		memory[16'h7698] <= 8'ha8;
		memory[16'h7699] <= 8'h42;
		memory[16'h769a] <= 8'h9e;
		memory[16'h769b] <= 8'ha5;
		memory[16'h769c] <= 8'h48;
		memory[16'h769d] <= 8'he7;
		memory[16'h769e] <= 8'h90;
		memory[16'h769f] <= 8'he2;
		memory[16'h76a0] <= 8'hc9;
		memory[16'h76a1] <= 8'hcf;
		memory[16'h76a2] <= 8'h72;
		memory[16'h76a3] <= 8'h86;
		memory[16'h76a4] <= 8'hae;
		memory[16'h76a5] <= 8'h24;
		memory[16'h76a6] <= 8'hd9;
		memory[16'h76a7] <= 8'he;
		memory[16'h76a8] <= 8'h5b;
		memory[16'h76a9] <= 8'hdb;
		memory[16'h76aa] <= 8'h72;
		memory[16'h76ab] <= 8'hb8;
		memory[16'h76ac] <= 8'h6c;
		memory[16'h76ad] <= 8'hd8;
		memory[16'h76ae] <= 8'h34;
		memory[16'h76af] <= 8'h45;
		memory[16'h76b0] <= 8'h85;
		memory[16'h76b1] <= 8'h74;
		memory[16'h76b2] <= 8'h4b;
		memory[16'h76b3] <= 8'hc6;
		memory[16'h76b4] <= 8'h7d;
		memory[16'h76b5] <= 8'hd2;
		memory[16'h76b6] <= 8'h15;
		memory[16'h76b7] <= 8'h25;
		memory[16'h76b8] <= 8'h15;
		memory[16'h76b9] <= 8'hb3;
		memory[16'h76ba] <= 8'hca;
		memory[16'h76bb] <= 8'h5d;
		memory[16'h76bc] <= 8'h9a;
		memory[16'h76bd] <= 8'h5b;
		memory[16'h76be] <= 8'h40;
		memory[16'h76bf] <= 8'h63;
		memory[16'h76c0] <= 8'h2a;
		memory[16'h76c1] <= 8'hb2;
		memory[16'h76c2] <= 8'he9;
		memory[16'h76c3] <= 8'hd8;
		memory[16'h76c4] <= 8'hd6;
		memory[16'h76c5] <= 8'hc3;
		memory[16'h76c6] <= 8'he6;
		memory[16'h76c7] <= 8'h31;
		memory[16'h76c8] <= 8'h9e;
		memory[16'h76c9] <= 8'h58;
		memory[16'h76ca] <= 8'he9;
		memory[16'h76cb] <= 8'ha;
		memory[16'h76cc] <= 8'h31;
		memory[16'h76cd] <= 8'h1d;
		memory[16'h76ce] <= 8'h4f;
		memory[16'h76cf] <= 8'hb6;
		memory[16'h76d0] <= 8'h92;
		memory[16'h76d1] <= 8'h9b;
		memory[16'h76d2] <= 8'h7c;
		memory[16'h76d3] <= 8'hf;
		memory[16'h76d4] <= 8'h6d;
		memory[16'h76d5] <= 8'h91;
		memory[16'h76d6] <= 8'h34;
		memory[16'h76d7] <= 8'h82;
		memory[16'h76d8] <= 8'h44;
		memory[16'h76d9] <= 8'hfe;
		memory[16'h76da] <= 8'he0;
		memory[16'h76db] <= 8'hde;
		memory[16'h76dc] <= 8'h59;
		memory[16'h76dd] <= 8'h20;
		memory[16'h76de] <= 8'h41;
		memory[16'h76df] <= 8'h83;
		memory[16'h76e0] <= 8'hd2;
		memory[16'h76e1] <= 8'h2a;
		memory[16'h76e2] <= 8'h5b;
		memory[16'h76e3] <= 8'ha8;
		memory[16'h76e4] <= 8'hed;
		memory[16'h76e5] <= 8'h41;
		memory[16'h76e6] <= 8'hd9;
		memory[16'h76e7] <= 8'h8b;
		memory[16'h76e8] <= 8'h9a;
		memory[16'h76e9] <= 8'hc2;
		memory[16'h76ea] <= 8'h95;
		memory[16'h76eb] <= 8'hcb;
		memory[16'h76ec] <= 8'hdf;
		memory[16'h76ed] <= 8'he5;
		memory[16'h76ee] <= 8'h81;
		memory[16'h76ef] <= 8'h71;
		memory[16'h76f0] <= 8'h80;
		memory[16'h76f1] <= 8'hfd;
		memory[16'h76f2] <= 8'h80;
		memory[16'h76f3] <= 8'hed;
		memory[16'h76f4] <= 8'h8e;
		memory[16'h76f5] <= 8'hb4;
		memory[16'h76f6] <= 8'h70;
		memory[16'h76f7] <= 8'hd2;
		memory[16'h76f8] <= 8'hb3;
		memory[16'h76f9] <= 8'h50;
		memory[16'h76fa] <= 8'hb0;
		memory[16'h76fb] <= 8'hc;
		memory[16'h76fc] <= 8'h70;
		memory[16'h76fd] <= 8'hf1;
		memory[16'h76fe] <= 8'h90;
		memory[16'h76ff] <= 8'h42;
		memory[16'h7700] <= 8'h1b;
		memory[16'h7701] <= 8'heb;
		memory[16'h7702] <= 8'hea;
		memory[16'h7703] <= 8'h9;
		memory[16'h7704] <= 8'h2d;
		memory[16'h7705] <= 8'hc3;
		memory[16'h7706] <= 8'h94;
		memory[16'h7707] <= 8'hc7;
		memory[16'h7708] <= 8'h85;
		memory[16'h7709] <= 8'h2a;
		memory[16'h770a] <= 8'h92;
		memory[16'h770b] <= 8'h64;
		memory[16'h770c] <= 8'hf;
		memory[16'h770d] <= 8'h13;
		memory[16'h770e] <= 8'hd6;
		memory[16'h770f] <= 8'h8f;
		memory[16'h7710] <= 8'h10;
		memory[16'h7711] <= 8'h56;
		memory[16'h7712] <= 8'h7c;
		memory[16'h7713] <= 8'h9e;
		memory[16'h7714] <= 8'hb;
		memory[16'h7715] <= 8'hec;
		memory[16'h7716] <= 8'h70;
		memory[16'h7717] <= 8'hbe;
		memory[16'h7718] <= 8'h3c;
		memory[16'h7719] <= 8'h20;
		memory[16'h771a] <= 8'hca;
		memory[16'h771b] <= 8'hac;
		memory[16'h771c] <= 8'h11;
		memory[16'h771d] <= 8'h5a;
		memory[16'h771e] <= 8'hee;
		memory[16'h771f] <= 8'h2c;
		memory[16'h7720] <= 8'h46;
		memory[16'h7721] <= 8'hd8;
		memory[16'h7722] <= 8'h35;
		memory[16'h7723] <= 8'h73;
		memory[16'h7724] <= 8'h9b;
		memory[16'h7725] <= 8'hca;
		memory[16'h7726] <= 8'h3a;
		memory[16'h7727] <= 8'h20;
		memory[16'h7728] <= 8'hf4;
		memory[16'h7729] <= 8'hcc;
		memory[16'h772a] <= 8'h85;
		memory[16'h772b] <= 8'h3;
		memory[16'h772c] <= 8'hdf;
		memory[16'h772d] <= 8'h5b;
		memory[16'h772e] <= 8'h92;
		memory[16'h772f] <= 8'hef;
		memory[16'h7730] <= 8'hb1;
		memory[16'h7731] <= 8'he;
		memory[16'h7732] <= 8'h8d;
		memory[16'h7733] <= 8'hbc;
		memory[16'h7734] <= 8'hfb;
		memory[16'h7735] <= 8'hfd;
		memory[16'h7736] <= 8'h7a;
		memory[16'h7737] <= 8'h37;
		memory[16'h7738] <= 8'h1d;
		memory[16'h7739] <= 8'h45;
		memory[16'h773a] <= 8'he4;
		memory[16'h773b] <= 8'h2e;
		memory[16'h773c] <= 8'h9f;
		memory[16'h773d] <= 8'hd2;
		memory[16'h773e] <= 8'h5a;
		memory[16'h773f] <= 8'he5;
		memory[16'h7740] <= 8'hab;
		memory[16'h7741] <= 8'h90;
		memory[16'h7742] <= 8'h58;
		memory[16'h7743] <= 8'h46;
		memory[16'h7744] <= 8'h5a;
		memory[16'h7745] <= 8'h92;
		memory[16'h7746] <= 8'h67;
		memory[16'h7747] <= 8'h4e;
		memory[16'h7748] <= 8'h5e;
		memory[16'h7749] <= 8'hec;
		memory[16'h774a] <= 8'h51;
		memory[16'h774b] <= 8'h3d;
		memory[16'h774c] <= 8'h47;
		memory[16'h774d] <= 8'he3;
		memory[16'h774e] <= 8'h2c;
		memory[16'h774f] <= 8'hf8;
		memory[16'h7750] <= 8'hf1;
		memory[16'h7751] <= 8'hb9;
		memory[16'h7752] <= 8'hb5;
		memory[16'h7753] <= 8'hec;
		memory[16'h7754] <= 8'hb6;
		memory[16'h7755] <= 8'h2f;
		memory[16'h7756] <= 8'h24;
		memory[16'h7757] <= 8'hd3;
		memory[16'h7758] <= 8'h74;
		memory[16'h7759] <= 8'h8;
		memory[16'h775a] <= 8'h1;
		memory[16'h775b] <= 8'h14;
		memory[16'h775c] <= 8'hda;
		memory[16'h775d] <= 8'h5c;
		memory[16'h775e] <= 8'hf9;
		memory[16'h775f] <= 8'h85;
		memory[16'h7760] <= 8'hec;
		memory[16'h7761] <= 8'h52;
		memory[16'h7762] <= 8'hcc;
		memory[16'h7763] <= 8'h46;
		memory[16'h7764] <= 8'he4;
		memory[16'h7765] <= 8'h33;
		memory[16'h7766] <= 8'h94;
		memory[16'h7767] <= 8'h43;
		memory[16'h7768] <= 8'h1f;
		memory[16'h7769] <= 8'he5;
		memory[16'h776a] <= 8'h80;
		memory[16'h776b] <= 8'h66;
		memory[16'h776c] <= 8'hc8;
		memory[16'h776d] <= 8'had;
		memory[16'h776e] <= 8'h5e;
		memory[16'h776f] <= 8'hb9;
		memory[16'h7770] <= 8'h66;
		memory[16'h7771] <= 8'h13;
		memory[16'h7772] <= 8'ha6;
		memory[16'h7773] <= 8'h1d;
		memory[16'h7774] <= 8'h43;
		memory[16'h7775] <= 8'hca;
		memory[16'h7776] <= 8'hf0;
		memory[16'h7777] <= 8'hb7;
		memory[16'h7778] <= 8'hd2;
		memory[16'h7779] <= 8'hf2;
		memory[16'h777a] <= 8'hcb;
		memory[16'h777b] <= 8'hac;
		memory[16'h777c] <= 8'h4e;
		memory[16'h777d] <= 8'hc5;
		memory[16'h777e] <= 8'h32;
		memory[16'h777f] <= 8'h3a;
		memory[16'h7780] <= 8'h17;
		memory[16'h7781] <= 8'hfe;
		memory[16'h7782] <= 8'h80;
		memory[16'h7783] <= 8'hfb;
		memory[16'h7784] <= 8'h31;
		memory[16'h7785] <= 8'h14;
		memory[16'h7786] <= 8'h3e;
		memory[16'h7787] <= 8'h50;
		memory[16'h7788] <= 8'hf9;
		memory[16'h7789] <= 8'hbf;
		memory[16'h778a] <= 8'hb6;
		memory[16'h778b] <= 8'hc1;
		memory[16'h778c] <= 8'h6c;
		memory[16'h778d] <= 8'h14;
		memory[16'h778e] <= 8'h7a;
		memory[16'h778f] <= 8'hd2;
		memory[16'h7790] <= 8'h28;
		memory[16'h7791] <= 8'h20;
		memory[16'h7792] <= 8'hef;
		memory[16'h7793] <= 8'h6b;
		memory[16'h7794] <= 8'hea;
		memory[16'h7795] <= 8'he0;
		memory[16'h7796] <= 8'h22;
		memory[16'h7797] <= 8'hbc;
		memory[16'h7798] <= 8'hd2;
		memory[16'h7799] <= 8'hee;
		memory[16'h779a] <= 8'h69;
		memory[16'h779b] <= 8'h20;
		memory[16'h779c] <= 8'hb3;
		memory[16'h779d] <= 8'h9b;
		memory[16'h779e] <= 8'h5a;
		memory[16'h779f] <= 8'hca;
		memory[16'h77a0] <= 8'h99;
		memory[16'h77a1] <= 8'hda;
		memory[16'h77a2] <= 8'hc5;
		memory[16'h77a3] <= 8'hca;
		memory[16'h77a4] <= 8'hee;
		memory[16'h77a5] <= 8'h4;
		memory[16'h77a6] <= 8'h1a;
		memory[16'h77a7] <= 8'he7;
		memory[16'h77a8] <= 8'hc3;
		memory[16'h77a9] <= 8'hd0;
		memory[16'h77aa] <= 8'ha8;
		memory[16'h77ab] <= 8'h2f;
		memory[16'h77ac] <= 8'he4;
		memory[16'h77ad] <= 8'h22;
		memory[16'h77ae] <= 8'h1;
		memory[16'h77af] <= 8'hc;
		memory[16'h77b0] <= 8'h43;
		memory[16'h77b1] <= 8'hf1;
		memory[16'h77b2] <= 8'h77;
		memory[16'h77b3] <= 8'h2d;
		memory[16'h77b4] <= 8'hd1;
		memory[16'h77b5] <= 8'h9a;
		memory[16'h77b6] <= 8'hea;
		memory[16'h77b7] <= 8'ha3;
		memory[16'h77b8] <= 8'h88;
		memory[16'h77b9] <= 8'h53;
		memory[16'h77ba] <= 8'hc3;
		memory[16'h77bb] <= 8'h3b;
		memory[16'h77bc] <= 8'hee;
		memory[16'h77bd] <= 8'h1d;
		memory[16'h77be] <= 8'h5;
		memory[16'h77bf] <= 8'h87;
		memory[16'h77c0] <= 8'hf7;
		memory[16'h77c1] <= 8'hca;
		memory[16'h77c2] <= 8'h51;
		memory[16'h77c3] <= 8'he5;
		memory[16'h77c4] <= 8'hce;
		memory[16'h77c5] <= 8'h6b;
		memory[16'h77c6] <= 8'hcc;
		memory[16'h77c7] <= 8'h91;
		memory[16'h77c8] <= 8'h3b;
		memory[16'h77c9] <= 8'h74;
		memory[16'h77ca] <= 8'hc0;
		memory[16'h77cb] <= 8'h1f;
		memory[16'h77cc] <= 8'h96;
		memory[16'h77cd] <= 8'hc2;
		memory[16'h77ce] <= 8'h2c;
		memory[16'h77cf] <= 8'hd9;
		memory[16'h77d0] <= 8'hb3;
		memory[16'h77d1] <= 8'ha3;
		memory[16'h77d2] <= 8'h7;
		memory[16'h77d3] <= 8'h84;
		memory[16'h77d4] <= 8'h3d;
		memory[16'h77d5] <= 8'hf1;
		memory[16'h77d6] <= 8'h27;
		memory[16'h77d7] <= 8'hc5;
		memory[16'h77d8] <= 8'h44;
		memory[16'h77d9] <= 8'hea;
		memory[16'h77da] <= 8'h0;
		memory[16'h77db] <= 8'h32;
		memory[16'h77dc] <= 8'h7;
		memory[16'h77dd] <= 8'h5;
		memory[16'h77de] <= 8'hb9;
		memory[16'h77df] <= 8'hfe;
		memory[16'h77e0] <= 8'hd0;
		memory[16'h77e1] <= 8'ha;
		memory[16'h77e2] <= 8'he3;
		memory[16'h77e3] <= 8'h9e;
		memory[16'h77e4] <= 8'h75;
		memory[16'h77e5] <= 8'haf;
		memory[16'h77e6] <= 8'h30;
		memory[16'h77e7] <= 8'hb0;
		memory[16'h77e8] <= 8'h23;
		memory[16'h77e9] <= 8'hf0;
		memory[16'h77ea] <= 8'hcf;
		memory[16'h77eb] <= 8'hb9;
		memory[16'h77ec] <= 8'hb2;
		memory[16'h77ed] <= 8'hfb;
		memory[16'h77ee] <= 8'h93;
		memory[16'h77ef] <= 8'h65;
		memory[16'h77f0] <= 8'h9f;
		memory[16'h77f1] <= 8'h9a;
		memory[16'h77f2] <= 8'he9;
		memory[16'h77f3] <= 8'hdc;
		memory[16'h77f4] <= 8'h8b;
		memory[16'h77f5] <= 8'h10;
		memory[16'h77f6] <= 8'ha2;
		memory[16'h77f7] <= 8'hcf;
		memory[16'h77f8] <= 8'hfa;
		memory[16'h77f9] <= 8'ha2;
		memory[16'h77fa] <= 8'h1;
		memory[16'h77fb] <= 8'h1;
		memory[16'h77fc] <= 8'ha8;
		memory[16'h77fd] <= 8'hba;
		memory[16'h77fe] <= 8'hff;
		memory[16'h77ff] <= 8'h78;
		memory[16'h7800] <= 8'hc4;
		memory[16'h7801] <= 8'he2;
		memory[16'h7802] <= 8'h16;
		memory[16'h7803] <= 8'h39;
		memory[16'h7804] <= 8'h91;
		memory[16'h7805] <= 8'h46;
		memory[16'h7806] <= 8'he9;
		memory[16'h7807] <= 8'hb4;
		memory[16'h7808] <= 8'h37;
		memory[16'h7809] <= 8'hb8;
		memory[16'h780a] <= 8'h6e;
		memory[16'h780b] <= 8'he9;
		memory[16'h780c] <= 8'hb4;
		memory[16'h780d] <= 8'h1;
		memory[16'h780e] <= 8'h4f;
		memory[16'h780f] <= 8'h53;
		memory[16'h7810] <= 8'h9b;
		memory[16'h7811] <= 8'h38;
		memory[16'h7812] <= 8'h2f;
		memory[16'h7813] <= 8'h26;
		memory[16'h7814] <= 8'h49;
		memory[16'h7815] <= 8'hd1;
		memory[16'h7816] <= 8'hf5;
		memory[16'h7817] <= 8'h43;
		memory[16'h7818] <= 8'h74;
		memory[16'h7819] <= 8'hf6;
		memory[16'h781a] <= 8'h45;
		memory[16'h781b] <= 8'h1c;
		memory[16'h781c] <= 8'hb0;
		memory[16'h781d] <= 8'h44;
		memory[16'h781e] <= 8'h94;
		memory[16'h781f] <= 8'h74;
		memory[16'h7820] <= 8'h27;
		memory[16'h7821] <= 8'haa;
		memory[16'h7822] <= 8'had;
		memory[16'h7823] <= 8'hb8;
		memory[16'h7824] <= 8'hf1;
		memory[16'h7825] <= 8'h96;
		memory[16'h7826] <= 8'h6d;
		memory[16'h7827] <= 8'h28;
		memory[16'h7828] <= 8'h4e;
		memory[16'h7829] <= 8'hdb;
		memory[16'h782a] <= 8'h11;
		memory[16'h782b] <= 8'h2;
		memory[16'h782c] <= 8'hdc;
		memory[16'h782d] <= 8'h60;
		memory[16'h782e] <= 8'h55;
		memory[16'h782f] <= 8'h77;
		memory[16'h7830] <= 8'h99;
		memory[16'h7831] <= 8'h85;
		memory[16'h7832] <= 8'h9d;
		memory[16'h7833] <= 8'he2;
		memory[16'h7834] <= 8'h56;
		memory[16'h7835] <= 8'h92;
		memory[16'h7836] <= 8'h25;
		memory[16'h7837] <= 8'hca;
		memory[16'h7838] <= 8'h88;
		memory[16'h7839] <= 8'h6a;
		memory[16'h783a] <= 8'he6;
		memory[16'h783b] <= 8'h38;
		memory[16'h783c] <= 8'haf;
		memory[16'h783d] <= 8'h7a;
		memory[16'h783e] <= 8'hac;
		memory[16'h783f] <= 8'hd6;
		memory[16'h7840] <= 8'h25;
		memory[16'h7841] <= 8'h59;
		memory[16'h7842] <= 8'h8e;
		memory[16'h7843] <= 8'h16;
		memory[16'h7844] <= 8'hef;
		memory[16'h7845] <= 8'hfb;
		memory[16'h7846] <= 8'h3e;
		memory[16'h7847] <= 8'h3d;
		memory[16'h7848] <= 8'hd6;
		memory[16'h7849] <= 8'h4f;
		memory[16'h784a] <= 8'h40;
		memory[16'h784b] <= 8'hb2;
		memory[16'h784c] <= 8'hb0;
		memory[16'h784d] <= 8'h95;
		memory[16'h784e] <= 8'h29;
		memory[16'h784f] <= 8'h49;
		memory[16'h7850] <= 8'h1a;
		memory[16'h7851] <= 8'hc6;
		memory[16'h7852] <= 8'h2b;
		memory[16'h7853] <= 8'h71;
		memory[16'h7854] <= 8'h58;
		memory[16'h7855] <= 8'h50;
		memory[16'h7856] <= 8'h3b;
		memory[16'h7857] <= 8'he0;
		memory[16'h7858] <= 8'hbb;
		memory[16'h7859] <= 8'h22;
		memory[16'h785a] <= 8'h18;
		memory[16'h785b] <= 8'h6a;
		memory[16'h785c] <= 8'h9c;
		memory[16'h785d] <= 8'hc4;
		memory[16'h785e] <= 8'h40;
		memory[16'h785f] <= 8'hc1;
		memory[16'h7860] <= 8'h1d;
		memory[16'h7861] <= 8'hce;
		memory[16'h7862] <= 8'hd7;
		memory[16'h7863] <= 8'hc;
		memory[16'h7864] <= 8'hca;
		memory[16'h7865] <= 8'h15;
		memory[16'h7866] <= 8'h4a;
		memory[16'h7867] <= 8'ha0;
		memory[16'h7868] <= 8'h65;
		memory[16'h7869] <= 8'h8a;
		memory[16'h786a] <= 8'h53;
		memory[16'h786b] <= 8'h15;
		memory[16'h786c] <= 8'h1f;
		memory[16'h786d] <= 8'h7c;
		memory[16'h786e] <= 8'h5e;
		memory[16'h786f] <= 8'h3a;
		memory[16'h7870] <= 8'h43;
		memory[16'h7871] <= 8'h89;
		memory[16'h7872] <= 8'hab;
		memory[16'h7873] <= 8'h9b;
		memory[16'h7874] <= 8'hd9;
		memory[16'h7875] <= 8'he6;
		memory[16'h7876] <= 8'h7c;
		memory[16'h7877] <= 8'h94;
		memory[16'h7878] <= 8'h8;
		memory[16'h7879] <= 8'h94;
		memory[16'h787a] <= 8'hfe;
		memory[16'h787b] <= 8'ha5;
		memory[16'h787c] <= 8'h59;
		memory[16'h787d] <= 8'h3e;
		memory[16'h787e] <= 8'h66;
		memory[16'h787f] <= 8'h76;
		memory[16'h7880] <= 8'hd;
		memory[16'h7881] <= 8'h3e;
		memory[16'h7882] <= 8'h83;
		memory[16'h7883] <= 8'hd7;
		memory[16'h7884] <= 8'h53;
		memory[16'h7885] <= 8'hcd;
		memory[16'h7886] <= 8'h77;
		memory[16'h7887] <= 8'hb8;
		memory[16'h7888] <= 8'h57;
		memory[16'h7889] <= 8'hca;
		memory[16'h788a] <= 8'hcd;
		memory[16'h788b] <= 8'h76;
		memory[16'h788c] <= 8'h47;
		memory[16'h788d] <= 8'h2b;
		memory[16'h788e] <= 8'hb0;
		memory[16'h788f] <= 8'h8a;
		memory[16'h7890] <= 8'hb4;
		memory[16'h7891] <= 8'h5b;
		memory[16'h7892] <= 8'h25;
		memory[16'h7893] <= 8'h8e;
		memory[16'h7894] <= 8'h42;
		memory[16'h7895] <= 8'ha1;
		memory[16'h7896] <= 8'h22;
		memory[16'h7897] <= 8'h4a;
		memory[16'h7898] <= 8'h36;
		memory[16'h7899] <= 8'h21;
		memory[16'h789a] <= 8'hef;
		memory[16'h789b] <= 8'h8f;
		memory[16'h789c] <= 8'h5f;
		memory[16'h789d] <= 8'h56;
		memory[16'h789e] <= 8'h5;
		memory[16'h789f] <= 8'h6c;
		memory[16'h78a0] <= 8'h94;
		memory[16'h78a1] <= 8'h88;
		memory[16'h78a2] <= 8'h43;
		memory[16'h78a3] <= 8'he7;
		memory[16'h78a4] <= 8'h55;
		memory[16'h78a5] <= 8'hbb;
		memory[16'h78a6] <= 8'ha0;
		memory[16'h78a7] <= 8'hac;
		memory[16'h78a8] <= 8'h85;
		memory[16'h78a9] <= 8'h6d;
		memory[16'h78aa] <= 8'h23;
		memory[16'h78ab] <= 8'hcc;
		memory[16'h78ac] <= 8'h99;
		memory[16'h78ad] <= 8'hd3;
		memory[16'h78ae] <= 8'h56;
		memory[16'h78af] <= 8'h4d;
		memory[16'h78b0] <= 8'h2f;
		memory[16'h78b1] <= 8'h7c;
		memory[16'h78b2] <= 8'hdb;
		memory[16'h78b3] <= 8'h71;
		memory[16'h78b4] <= 8'h1d;
		memory[16'h78b5] <= 8'hfe;
		memory[16'h78b6] <= 8'hbb;
		memory[16'h78b7] <= 8'h53;
		memory[16'h78b8] <= 8'h1f;
		memory[16'h78b9] <= 8'hab;
		memory[16'h78ba] <= 8'he2;
		memory[16'h78bb] <= 8'h7e;
		memory[16'h78bc] <= 8'h1;
		memory[16'h78bd] <= 8'he8;
		memory[16'h78be] <= 8'heb;
		memory[16'h78bf] <= 8'h95;
		memory[16'h78c0] <= 8'h70;
		memory[16'h78c1] <= 8'h2e;
		memory[16'h78c2] <= 8'h7c;
		memory[16'h78c3] <= 8'hc6;
		memory[16'h78c4] <= 8'he9;
		memory[16'h78c5] <= 8'h1c;
		memory[16'h78c6] <= 8'h72;
		memory[16'h78c7] <= 8'h6f;
		memory[16'h78c8] <= 8'h8a;
		memory[16'h78c9] <= 8'h95;
		memory[16'h78ca] <= 8'h3b;
		memory[16'h78cb] <= 8'h23;
		memory[16'h78cc] <= 8'h69;
		memory[16'h78cd] <= 8'h92;
		memory[16'h78ce] <= 8'h70;
		memory[16'h78cf] <= 8'h98;
		memory[16'h78d0] <= 8'he;
		memory[16'h78d1] <= 8'h4c;
		memory[16'h78d2] <= 8'h9;
		memory[16'h78d3] <= 8'h2b;
		memory[16'h78d4] <= 8'h4a;
		memory[16'h78d5] <= 8'hc4;
		memory[16'h78d6] <= 8'h7f;
		memory[16'h78d7] <= 8'h69;
		memory[16'h78d8] <= 8'h6f;
		memory[16'h78d9] <= 8'h61;
		memory[16'h78da] <= 8'he7;
		memory[16'h78db] <= 8'h70;
		memory[16'h78dc] <= 8'h49;
		memory[16'h78dd] <= 8'hd2;
		memory[16'h78de] <= 8'h5;
		memory[16'h78df] <= 8'hba;
		memory[16'h78e0] <= 8'h1;
		memory[16'h78e1] <= 8'h82;
		memory[16'h78e2] <= 8'h80;
		memory[16'h78e3] <= 8'hea;
		memory[16'h78e4] <= 8'h9e;
		memory[16'h78e5] <= 8'hf2;
		memory[16'h78e6] <= 8'h59;
		memory[16'h78e7] <= 8'h28;
		memory[16'h78e8] <= 8'h88;
		memory[16'h78e9] <= 8'h95;
		memory[16'h78ea] <= 8'h4b;
		memory[16'h78eb] <= 8'hf1;
		memory[16'h78ec] <= 8'h27;
		memory[16'h78ed] <= 8'hbc;
		memory[16'h78ee] <= 8'h89;
		memory[16'h78ef] <= 8'h35;
		memory[16'h78f0] <= 8'h8;
		memory[16'h78f1] <= 8'h92;
		memory[16'h78f2] <= 8'h60;
		memory[16'h78f3] <= 8'h52;
		memory[16'h78f4] <= 8'h56;
		memory[16'h78f5] <= 8'hdf;
		memory[16'h78f6] <= 8'hbb;
		memory[16'h78f7] <= 8'hc6;
		memory[16'h78f8] <= 8'h41;
		memory[16'h78f9] <= 8'ha2;
		memory[16'h78fa] <= 8'h36;
		memory[16'h78fb] <= 8'h8a;
		memory[16'h78fc] <= 8'h75;
		memory[16'h78fd] <= 8'h3c;
		memory[16'h78fe] <= 8'h44;
		memory[16'h78ff] <= 8'h76;
		memory[16'h7900] <= 8'hbe;
		memory[16'h7901] <= 8'hc4;
		memory[16'h7902] <= 8'h60;
		memory[16'h7903] <= 8'h5c;
		memory[16'h7904] <= 8'hb7;
		memory[16'h7905] <= 8'hba;
		memory[16'h7906] <= 8'h85;
		memory[16'h7907] <= 8'h3f;
		memory[16'h7908] <= 8'h4f;
		memory[16'h7909] <= 8'hd0;
		memory[16'h790a] <= 8'h30;
		memory[16'h790b] <= 8'h76;
		memory[16'h790c] <= 8'h8c;
		memory[16'h790d] <= 8'hb9;
		memory[16'h790e] <= 8'hab;
		memory[16'h790f] <= 8'h94;
		memory[16'h7910] <= 8'h4b;
		memory[16'h7911] <= 8'hb;
		memory[16'h7912] <= 8'he6;
		memory[16'h7913] <= 8'ha1;
		memory[16'h7914] <= 8'heb;
		memory[16'h7915] <= 8'ha1;
		memory[16'h7916] <= 8'h67;
		memory[16'h7917] <= 8'h2c;
		memory[16'h7918] <= 8'h44;
		memory[16'h7919] <= 8'h9e;
		memory[16'h791a] <= 8'hb6;
		memory[16'h791b] <= 8'hb9;
		memory[16'h791c] <= 8'hda;
		memory[16'h791d] <= 8'hfb;
		memory[16'h791e] <= 8'h2f;
		memory[16'h791f] <= 8'h98;
		memory[16'h7920] <= 8'hbf;
		memory[16'h7921] <= 8'h8f;
		memory[16'h7922] <= 8'hf4;
		memory[16'h7923] <= 8'h76;
		memory[16'h7924] <= 8'h49;
		memory[16'h7925] <= 8'h79;
		memory[16'h7926] <= 8'hb5;
		memory[16'h7927] <= 8'h98;
		memory[16'h7928] <= 8'h4a;
		memory[16'h7929] <= 8'he5;
		memory[16'h792a] <= 8'he;
		memory[16'h792b] <= 8'hd6;
		memory[16'h792c] <= 8'h9e;
		memory[16'h792d] <= 8'hb9;
		memory[16'h792e] <= 8'h6b;
		memory[16'h792f] <= 8'he9;
		memory[16'h7930] <= 8'hc5;
		memory[16'h7931] <= 8'h51;
		memory[16'h7932] <= 8'h8b;
		memory[16'h7933] <= 8'hb0;
		memory[16'h7934] <= 8'hf3;
		memory[16'h7935] <= 8'hf2;
		memory[16'h7936] <= 8'hdc;
		memory[16'h7937] <= 8'h37;
		memory[16'h7938] <= 8'h90;
		memory[16'h7939] <= 8'h92;
		memory[16'h793a] <= 8'hf0;
		memory[16'h793b] <= 8'h6a;
		memory[16'h793c] <= 8'h8d;
		memory[16'h793d] <= 8'h1f;
		memory[16'h793e] <= 8'h2;
		memory[16'h793f] <= 8'h4d;
		memory[16'h7940] <= 8'hae;
		memory[16'h7941] <= 8'hf7;
		memory[16'h7942] <= 8'hc3;
		memory[16'h7943] <= 8'hf8;
		memory[16'h7944] <= 8'h70;
		memory[16'h7945] <= 8'h79;
		memory[16'h7946] <= 8'h90;
		memory[16'h7947] <= 8'hba;
		memory[16'h7948] <= 8'h5e;
		memory[16'h7949] <= 8'h9f;
		memory[16'h794a] <= 8'h91;
		memory[16'h794b] <= 8'hfd;
		memory[16'h794c] <= 8'h58;
		memory[16'h794d] <= 8'hfc;
		memory[16'h794e] <= 8'he6;
		memory[16'h794f] <= 8'h1d;
		memory[16'h7950] <= 8'h4d;
		memory[16'h7951] <= 8'h71;
		memory[16'h7952] <= 8'hcd;
		memory[16'h7953] <= 8'h40;
		memory[16'h7954] <= 8'h64;
		memory[16'h7955] <= 8'ha9;
		memory[16'h7956] <= 8'h77;
		memory[16'h7957] <= 8'hf4;
		memory[16'h7958] <= 8'h3c;
		memory[16'h7959] <= 8'h67;
		memory[16'h795a] <= 8'h5f;
		memory[16'h795b] <= 8'hc9;
		memory[16'h795c] <= 8'h86;
		memory[16'h795d] <= 8'h61;
		memory[16'h795e] <= 8'h16;
		memory[16'h795f] <= 8'h35;
		memory[16'h7960] <= 8'h58;
		memory[16'h7961] <= 8'hda;
		memory[16'h7962] <= 8'h2d;
		memory[16'h7963] <= 8'hc9;
		memory[16'h7964] <= 8'h53;
		memory[16'h7965] <= 8'hbd;
		memory[16'h7966] <= 8'h83;
		memory[16'h7967] <= 8'hb1;
		memory[16'h7968] <= 8'h5c;
		memory[16'h7969] <= 8'h14;
		memory[16'h796a] <= 8'hae;
		memory[16'h796b] <= 8'hb5;
		memory[16'h796c] <= 8'h10;
		memory[16'h796d] <= 8'h95;
		memory[16'h796e] <= 8'hd2;
		memory[16'h796f] <= 8'h5e;
		memory[16'h7970] <= 8'h6;
		memory[16'h7971] <= 8'ha0;
		memory[16'h7972] <= 8'h9e;
		memory[16'h7973] <= 8'h6a;
		memory[16'h7974] <= 8'h49;
		memory[16'h7975] <= 8'h16;
		memory[16'h7976] <= 8'h5f;
		memory[16'h7977] <= 8'h85;
		memory[16'h7978] <= 8'h7d;
		memory[16'h7979] <= 8'hbe;
		memory[16'h797a] <= 8'h4f;
		memory[16'h797b] <= 8'h4;
		memory[16'h797c] <= 8'h1f;
		memory[16'h797d] <= 8'h65;
		memory[16'h797e] <= 8'h39;
		memory[16'h797f] <= 8'h78;
		memory[16'h7980] <= 8'h3f;
		memory[16'h7981] <= 8'h66;
		memory[16'h7982] <= 8'h41;
		memory[16'h7983] <= 8'h92;
		memory[16'h7984] <= 8'h23;
		memory[16'h7985] <= 8'hc4;
		memory[16'h7986] <= 8'h44;
		memory[16'h7987] <= 8'h80;
		memory[16'h7988] <= 8'hd9;
		memory[16'h7989] <= 8'hf2;
		memory[16'h798a] <= 8'h35;
		memory[16'h798b] <= 8'he9;
		memory[16'h798c] <= 8'h87;
		memory[16'h798d] <= 8'h7;
		memory[16'h798e] <= 8'h47;
		memory[16'h798f] <= 8'h8e;
		memory[16'h7990] <= 8'ha7;
		memory[16'h7991] <= 8'he6;
		memory[16'h7992] <= 8'hf8;
		memory[16'h7993] <= 8'hf1;
		memory[16'h7994] <= 8'hfc;
		memory[16'h7995] <= 8'h57;
		memory[16'h7996] <= 8'h76;
		memory[16'h7997] <= 8'h79;
		memory[16'h7998] <= 8'h15;
		memory[16'h7999] <= 8'hc5;
		memory[16'h799a] <= 8'h7d;
		memory[16'h799b] <= 8'h35;
		memory[16'h799c] <= 8'h2b;
		memory[16'h799d] <= 8'hb6;
		memory[16'h799e] <= 8'had;
		memory[16'h799f] <= 8'h6a;
		memory[16'h79a0] <= 8'h1c;
		memory[16'h79a1] <= 8'hee;
		memory[16'h79a2] <= 8'hfd;
		memory[16'h79a3] <= 8'h40;
		memory[16'h79a4] <= 8'hb2;
		memory[16'h79a5] <= 8'h41;
		memory[16'h79a6] <= 8'hc0;
		memory[16'h79a7] <= 8'h8b;
		memory[16'h79a8] <= 8'h33;
		memory[16'h79a9] <= 8'hf5;
		memory[16'h79aa] <= 8'h75;
		memory[16'h79ab] <= 8'hbb;
		memory[16'h79ac] <= 8'hfc;
		memory[16'h79ad] <= 8'hbc;
		memory[16'h79ae] <= 8'h49;
		memory[16'h79af] <= 8'ha4;
		memory[16'h79b0] <= 8'ha2;
		memory[16'h79b1] <= 8'h41;
		memory[16'h79b2] <= 8'h95;
		memory[16'h79b3] <= 8'h9e;
		memory[16'h79b4] <= 8'h99;
		memory[16'h79b5] <= 8'hb;
		memory[16'h79b6] <= 8'h18;
		memory[16'h79b7] <= 8'hae;
		memory[16'h79b8] <= 8'hd1;
		memory[16'h79b9] <= 8'h95;
		memory[16'h79ba] <= 8'he3;
		memory[16'h79bb] <= 8'hfc;
		memory[16'h79bc] <= 8'h4c;
		memory[16'h79bd] <= 8'h90;
		memory[16'h79be] <= 8'h66;
		memory[16'h79bf] <= 8'h68;
		memory[16'h79c0] <= 8'h7e;
		memory[16'h79c1] <= 8'h63;
		memory[16'h79c2] <= 8'ha8;
		memory[16'h79c3] <= 8'h31;
		memory[16'h79c4] <= 8'ha4;
		memory[16'h79c5] <= 8'h68;
		memory[16'h79c6] <= 8'hbc;
		memory[16'h79c7] <= 8'hd8;
		memory[16'h79c8] <= 8'h5d;
		memory[16'h79c9] <= 8'h31;
		memory[16'h79ca] <= 8'h93;
		memory[16'h79cb] <= 8'h5a;
		memory[16'h79cc] <= 8'hee;
		memory[16'h79cd] <= 8'hdc;
		memory[16'h79ce] <= 8'hfe;
		memory[16'h79cf] <= 8'h90;
		memory[16'h79d0] <= 8'h1d;
		memory[16'h79d1] <= 8'h93;
		memory[16'h79d2] <= 8'h2f;
		memory[16'h79d3] <= 8'hb6;
		memory[16'h79d4] <= 8'h9e;
		memory[16'h79d5] <= 8'h47;
		memory[16'h79d6] <= 8'h65;
		memory[16'h79d7] <= 8'h6f;
		memory[16'h79d8] <= 8'hdc;
		memory[16'h79d9] <= 8'h48;
		memory[16'h79da] <= 8'h6b;
		memory[16'h79db] <= 8'h28;
		memory[16'h79dc] <= 8'hd9;
		memory[16'h79dd] <= 8'hd2;
		memory[16'h79de] <= 8'h91;
		memory[16'h79df] <= 8'h57;
		memory[16'h79e0] <= 8'h35;
		memory[16'h79e1] <= 8'h39;
		memory[16'h79e2] <= 8'h88;
		memory[16'h79e3] <= 8'hda;
		memory[16'h79e4] <= 8'ha2;
		memory[16'h79e5] <= 8'h45;
		memory[16'h79e6] <= 8'hb2;
		memory[16'h79e7] <= 8'hff;
		memory[16'h79e8] <= 8'h76;
		memory[16'h79e9] <= 8'h45;
		memory[16'h79ea] <= 8'h59;
		memory[16'h79eb] <= 8'h64;
		memory[16'h79ec] <= 8'h21;
		memory[16'h79ed] <= 8'h57;
		memory[16'h79ee] <= 8'hf5;
		memory[16'h79ef] <= 8'h3e;
		memory[16'h79f0] <= 8'hea;
		memory[16'h79f1] <= 8'h24;
		memory[16'h79f2] <= 8'hf5;
		memory[16'h79f3] <= 8'h89;
		memory[16'h79f4] <= 8'h6b;
		memory[16'h79f5] <= 8'h5a;
		memory[16'h79f6] <= 8'hf8;
		memory[16'h79f7] <= 8'h47;
		memory[16'h79f8] <= 8'ha2;
		memory[16'h79f9] <= 8'h64;
		memory[16'h79fa] <= 8'h70;
		memory[16'h79fb] <= 8'h7b;
		memory[16'h79fc] <= 8'h36;
		memory[16'h79fd] <= 8'h1;
		memory[16'h79fe] <= 8'hd3;
		memory[16'h79ff] <= 8'h6b;
		memory[16'h7a00] <= 8'h3a;
		memory[16'h7a01] <= 8'h5b;
		memory[16'h7a02] <= 8'h45;
		memory[16'h7a03] <= 8'hdc;
		memory[16'h7a04] <= 8'ha0;
		memory[16'h7a05] <= 8'hf7;
		memory[16'h7a06] <= 8'hdc;
		memory[16'h7a07] <= 8'h17;
		memory[16'h7a08] <= 8'h3c;
		memory[16'h7a09] <= 8'h35;
		memory[16'h7a0a] <= 8'h7b;
		memory[16'h7a0b] <= 8'h5d;
		memory[16'h7a0c] <= 8'h8d;
		memory[16'h7a0d] <= 8'h70;
		memory[16'h7a0e] <= 8'h9c;
		memory[16'h7a0f] <= 8'h77;
		memory[16'h7a10] <= 8'h94;
		memory[16'h7a11] <= 8'h91;
		memory[16'h7a12] <= 8'h0;
		memory[16'h7a13] <= 8'hff;
		memory[16'h7a14] <= 8'heb;
		memory[16'h7a15] <= 8'hf9;
		memory[16'h7a16] <= 8'h47;
		memory[16'h7a17] <= 8'h8d;
		memory[16'h7a18] <= 8'h5d;
		memory[16'h7a19] <= 8'hb7;
		memory[16'h7a1a] <= 8'h9;
		memory[16'h7a1b] <= 8'h93;
		memory[16'h7a1c] <= 8'hb8;
		memory[16'h7a1d] <= 8'hdc;
		memory[16'h7a1e] <= 8'hfe;
		memory[16'h7a1f] <= 8'hf2;
		memory[16'h7a20] <= 8'h37;
		memory[16'h7a21] <= 8'h44;
		memory[16'h7a22] <= 8'hcf;
		memory[16'h7a23] <= 8'hd8;
		memory[16'h7a24] <= 8'h3b;
		memory[16'h7a25] <= 8'hab;
		memory[16'h7a26] <= 8'hef;
		memory[16'h7a27] <= 8'h78;
		memory[16'h7a28] <= 8'he0;
		memory[16'h7a29] <= 8'h6a;
		memory[16'h7a2a] <= 8'hd5;
		memory[16'h7a2b] <= 8'h6d;
		memory[16'h7a2c] <= 8'hdb;
		memory[16'h7a2d] <= 8'h71;
		memory[16'h7a2e] <= 8'he5;
		memory[16'h7a2f] <= 8'h6f;
		memory[16'h7a30] <= 8'h2;
		memory[16'h7a31] <= 8'he5;
		memory[16'h7a32] <= 8'h6f;
		memory[16'h7a33] <= 8'hed;
		memory[16'h7a34] <= 8'hde;
		memory[16'h7a35] <= 8'hb6;
		memory[16'h7a36] <= 8'h7b;
		memory[16'h7a37] <= 8'h3b;
		memory[16'h7a38] <= 8'h6d;
		memory[16'h7a39] <= 8'h84;
		memory[16'h7a3a] <= 8'hce;
		memory[16'h7a3b] <= 8'h25;
		memory[16'h7a3c] <= 8'h60;
		memory[16'h7a3d] <= 8'hcd;
		memory[16'h7a3e] <= 8'h17;
		memory[16'h7a3f] <= 8'h97;
		memory[16'h7a40] <= 8'h11;
		memory[16'h7a41] <= 8'he6;
		memory[16'h7a42] <= 8'h6f;
		memory[16'h7a43] <= 8'h4c;
		memory[16'h7a44] <= 8'h91;
		memory[16'h7a45] <= 8'h5e;
		memory[16'h7a46] <= 8'hc4;
		memory[16'h7a47] <= 8'h72;
		memory[16'h7a48] <= 8'hc9;
		memory[16'h7a49] <= 8'h9a;
		memory[16'h7a4a] <= 8'hdf;
		memory[16'h7a4b] <= 8'ha4;
		memory[16'h7a4c] <= 8'hb;
		memory[16'h7a4d] <= 8'hc4;
		memory[16'h7a4e] <= 8'h13;
		memory[16'h7a4f] <= 8'he;
		memory[16'h7a50] <= 8'haa;
		memory[16'h7a51] <= 8'h82;
		memory[16'h7a52] <= 8'hfb;
		memory[16'h7a53] <= 8'h88;
		memory[16'h7a54] <= 8'h38;
		memory[16'h7a55] <= 8'h76;
		memory[16'h7a56] <= 8'hc4;
		memory[16'h7a57] <= 8'ha5;
		memory[16'h7a58] <= 8'hfa;
		memory[16'h7a59] <= 8'h92;
		memory[16'h7a5a] <= 8'hca;
		memory[16'h7a5b] <= 8'h5a;
		memory[16'h7a5c] <= 8'h5f;
		memory[16'h7a5d] <= 8'he2;
		memory[16'h7a5e] <= 8'hf2;
		memory[16'h7a5f] <= 8'h70;
		memory[16'h7a60] <= 8'hc8;
		memory[16'h7a61] <= 8'h61;
		memory[16'h7a62] <= 8'hbd;
		memory[16'h7a63] <= 8'h5a;
		memory[16'h7a64] <= 8'hc0;
		memory[16'h7a65] <= 8'h81;
		memory[16'h7a66] <= 8'hcc;
		memory[16'h7a67] <= 8'h89;
		memory[16'h7a68] <= 8'h1b;
		memory[16'h7a69] <= 8'hab;
		memory[16'h7a6a] <= 8'h2d;
		memory[16'h7a6b] <= 8'h27;
		memory[16'h7a6c] <= 8'h70;
		memory[16'h7a6d] <= 8'h40;
		memory[16'h7a6e] <= 8'h35;
		memory[16'h7a6f] <= 8'h1a;
		memory[16'h7a70] <= 8'hc3;
		memory[16'h7a71] <= 8'h30;
		memory[16'h7a72] <= 8'ha2;
		memory[16'h7a73] <= 8'hfb;
		memory[16'h7a74] <= 8'ha7;
		memory[16'h7a75] <= 8'h66;
		memory[16'h7a76] <= 8'ha1;
		memory[16'h7a77] <= 8'ha1;
		memory[16'h7a78] <= 8'hf9;
		memory[16'h7a79] <= 8'h6b;
		memory[16'h7a7a] <= 8'hfc;
		memory[16'h7a7b] <= 8'h58;
		memory[16'h7a7c] <= 8'h4d;
		memory[16'h7a7d] <= 8'hee;
		memory[16'h7a7e] <= 8'hc9;
		memory[16'h7a7f] <= 8'h16;
		memory[16'h7a80] <= 8'h4f;
		memory[16'h7a81] <= 8'h86;
		memory[16'h7a82] <= 8'h70;
		memory[16'h7a83] <= 8'hf;
		memory[16'h7a84] <= 8'h7;
		memory[16'h7a85] <= 8'h3c;
		memory[16'h7a86] <= 8'h98;
		memory[16'h7a87] <= 8'h23;
		memory[16'h7a88] <= 8'he7;
		memory[16'h7a89] <= 8'hc5;
		memory[16'h7a8a] <= 8'h4a;
		memory[16'h7a8b] <= 8'h57;
		memory[16'h7a8c] <= 8'h6;
		memory[16'h7a8d] <= 8'h7f;
		memory[16'h7a8e] <= 8'h71;
		memory[16'h7a8f] <= 8'hc9;
		memory[16'h7a90] <= 8'haf;
		memory[16'h7a91] <= 8'h14;
		memory[16'h7a92] <= 8'hc4;
		memory[16'h7a93] <= 8'h56;
		memory[16'h7a94] <= 8'h7a;
		memory[16'h7a95] <= 8'h65;
		memory[16'h7a96] <= 8'hf8;
		memory[16'h7a97] <= 8'h73;
		memory[16'h7a98] <= 8'hd1;
		memory[16'h7a99] <= 8'hf4;
		memory[16'h7a9a] <= 8'hcc;
		memory[16'h7a9b] <= 8'h1e;
		memory[16'h7a9c] <= 8'he2;
		memory[16'h7a9d] <= 8'h95;
		memory[16'h7a9e] <= 8'h34;
		memory[16'h7a9f] <= 8'h31;
		memory[16'h7aa0] <= 8'h1b;
		memory[16'h7aa1] <= 8'ha4;
		memory[16'h7aa2] <= 8'h41;
		memory[16'h7aa3] <= 8'h22;
		memory[16'h7aa4] <= 8'he0;
		memory[16'h7aa5] <= 8'hd9;
		memory[16'h7aa6] <= 8'h45;
		memory[16'h7aa7] <= 8'hc8;
		memory[16'h7aa8] <= 8'h9f;
		memory[16'h7aa9] <= 8'h8f;
		memory[16'h7aaa] <= 8'h1f;
		memory[16'h7aab] <= 8'ha5;
		memory[16'h7aac] <= 8'he;
		memory[16'h7aad] <= 8'h91;
		memory[16'h7aae] <= 8'h6e;
		memory[16'h7aaf] <= 8'hbe;
		memory[16'h7ab0] <= 8'ha5;
		memory[16'h7ab1] <= 8'h32;
		memory[16'h7ab2] <= 8'h14;
		memory[16'h7ab3] <= 8'h1f;
		memory[16'h7ab4] <= 8'h98;
		memory[16'h7ab5] <= 8'hc;
		memory[16'h7ab6] <= 8'h93;
		memory[16'h7ab7] <= 8'h69;
		memory[16'h7ab8] <= 8'h0;
		memory[16'h7ab9] <= 8'h5f;
		memory[16'h7aba] <= 8'h87;
		memory[16'h7abb] <= 8'he2;
		memory[16'h7abc] <= 8'hf4;
		memory[16'h7abd] <= 8'hbc;
		memory[16'h7abe] <= 8'h14;
		memory[16'h7abf] <= 8'hf;
		memory[16'h7ac0] <= 8'h60;
		memory[16'h7ac1] <= 8'h55;
		memory[16'h7ac2] <= 8'h31;
		memory[16'h7ac3] <= 8'h41;
		memory[16'h7ac4] <= 8'h2e;
		memory[16'h7ac5] <= 8'h77;
		memory[16'h7ac6] <= 8'h9;
		memory[16'h7ac7] <= 8'hcd;
		memory[16'h7ac8] <= 8'h6;
		memory[16'h7ac9] <= 8'h28;
		memory[16'h7aca] <= 8'h72;
		memory[16'h7acb] <= 8'h15;
		memory[16'h7acc] <= 8'hb9;
		memory[16'h7acd] <= 8'he0;
		memory[16'h7ace] <= 8'hd3;
		memory[16'h7acf] <= 8'h5e;
		memory[16'h7ad0] <= 8'h13;
		memory[16'h7ad1] <= 8'he7;
		memory[16'h7ad2] <= 8'h7e;
		memory[16'h7ad3] <= 8'hab;
		memory[16'h7ad4] <= 8'hf4;
		memory[16'h7ad5] <= 8'h11;
		memory[16'h7ad6] <= 8'h14;
		memory[16'h7ad7] <= 8'hf4;
		memory[16'h7ad8] <= 8'h70;
		memory[16'h7ad9] <= 8'h9b;
		memory[16'h7ada] <= 8'hd7;
		memory[16'h7adb] <= 8'h64;
		memory[16'h7adc] <= 8'h57;
		memory[16'h7add] <= 8'heb;
		memory[16'h7ade] <= 8'h73;
		memory[16'h7adf] <= 8'hb8;
		memory[16'h7ae0] <= 8'h40;
		memory[16'h7ae1] <= 8'ha4;
		memory[16'h7ae2] <= 8'hf9;
		memory[16'h7ae3] <= 8'h6e;
		memory[16'h7ae4] <= 8'h1b;
		memory[16'h7ae5] <= 8'h2;
		memory[16'h7ae6] <= 8'h3c;
		memory[16'h7ae7] <= 8'h22;
		memory[16'h7ae8] <= 8'h2a;
		memory[16'h7ae9] <= 8'hae;
		memory[16'h7aea] <= 8'h37;
		memory[16'h7aeb] <= 8'he4;
		memory[16'h7aec] <= 8'h8f;
		memory[16'h7aed] <= 8'ha;
		memory[16'h7aee] <= 8'h42;
		memory[16'h7aef] <= 8'ha2;
		memory[16'h7af0] <= 8'hf1;
		memory[16'h7af1] <= 8'hc0;
		memory[16'h7af2] <= 8'h4d;
		memory[16'h7af3] <= 8'he5;
		memory[16'h7af4] <= 8'hd1;
		memory[16'h7af5] <= 8'h61;
		memory[16'h7af6] <= 8'hda;
		memory[16'h7af7] <= 8'h41;
		memory[16'h7af8] <= 8'hfc;
		memory[16'h7af9] <= 8'hb1;
		memory[16'h7afa] <= 8'ha5;
		memory[16'h7afb] <= 8'h54;
		memory[16'h7afc] <= 8'h9c;
		memory[16'h7afd] <= 8'h18;
		memory[16'h7afe] <= 8'hc;
		memory[16'h7aff] <= 8'hdc;
		memory[16'h7b00] <= 8'hbd;
		memory[16'h7b01] <= 8'h5;
		memory[16'h7b02] <= 8'h4a;
		memory[16'h7b03] <= 8'hd8;
		memory[16'h7b04] <= 8'h7;
		memory[16'h7b05] <= 8'h86;
		memory[16'h7b06] <= 8'hfa;
		memory[16'h7b07] <= 8'h31;
		memory[16'h7b08] <= 8'h35;
		memory[16'h7b09] <= 8'h31;
		memory[16'h7b0a] <= 8'h15;
		memory[16'h7b0b] <= 8'hc4;
		memory[16'h7b0c] <= 8'h3b;
		memory[16'h7b0d] <= 8'h58;
		memory[16'h7b0e] <= 8'h66;
		memory[16'h7b0f] <= 8'h2d;
		memory[16'h7b10] <= 8'h18;
		memory[16'h7b11] <= 8'hb3;
		memory[16'h7b12] <= 8'h12;
		memory[16'h7b13] <= 8'hea;
		memory[16'h7b14] <= 8'h14;
		memory[16'h7b15] <= 8'hec;
		memory[16'h7b16] <= 8'h2b;
		memory[16'h7b17] <= 8'h10;
		memory[16'h7b18] <= 8'h9d;
		memory[16'h7b19] <= 8'hd1;
		memory[16'h7b1a] <= 8'h64;
		memory[16'h7b1b] <= 8'h39;
		memory[16'h7b1c] <= 8'he9;
		memory[16'h7b1d] <= 8'h70;
		memory[16'h7b1e] <= 8'h15;
		memory[16'h7b1f] <= 8'ha6;
		memory[16'h7b20] <= 8'h75;
		memory[16'h7b21] <= 8'h60;
		memory[16'h7b22] <= 8'h7f;
		memory[16'h7b23] <= 8'h7c;
		memory[16'h7b24] <= 8'he6;
		memory[16'h7b25] <= 8'h79;
		memory[16'h7b26] <= 8'hae;
		memory[16'h7b27] <= 8'h1b;
		memory[16'h7b28] <= 8'hab;
		memory[16'h7b29] <= 8'hc3;
		memory[16'h7b2a] <= 8'hdf;
		memory[16'h7b2b] <= 8'he6;
		memory[16'h7b2c] <= 8'h1b;
		memory[16'h7b2d] <= 8'h45;
		memory[16'h7b2e] <= 8'h13;
		memory[16'h7b2f] <= 8'h34;
		memory[16'h7b30] <= 8'hf8;
		memory[16'h7b31] <= 8'h26;
		memory[16'h7b32] <= 8'h1e;
		memory[16'h7b33] <= 8'hc;
		memory[16'h7b34] <= 8'h12;
		memory[16'h7b35] <= 8'h49;
		memory[16'h7b36] <= 8'h1d;
		memory[16'h7b37] <= 8'hb0;
		memory[16'h7b38] <= 8'h1a;
		memory[16'h7b39] <= 8'h81;
		memory[16'h7b3a] <= 8'he9;
		memory[16'h7b3b] <= 8'h4;
		memory[16'h7b3c] <= 8'hf2;
		memory[16'h7b3d] <= 8'hff;
		memory[16'h7b3e] <= 8'haa;
		memory[16'h7b3f] <= 8'h67;
		memory[16'h7b40] <= 8'h5f;
		memory[16'h7b41] <= 8'h29;
		memory[16'h7b42] <= 8'he4;
		memory[16'h7b43] <= 8'h45;
		memory[16'h7b44] <= 8'ha3;
		memory[16'h7b45] <= 8'h92;
		memory[16'h7b46] <= 8'h61;
		memory[16'h7b47] <= 8'h4e;
		memory[16'h7b48] <= 8'h55;
		memory[16'h7b49] <= 8'h40;
		memory[16'h7b4a] <= 8'h34;
		memory[16'h7b4b] <= 8'h71;
		memory[16'h7b4c] <= 8'h86;
		memory[16'h7b4d] <= 8'h48;
		memory[16'h7b4e] <= 8'ha5;
		memory[16'h7b4f] <= 8'h7e;
		memory[16'h7b50] <= 8'h6e;
		memory[16'h7b51] <= 8'hc3;
		memory[16'h7b52] <= 8'h8b;
		memory[16'h7b53] <= 8'h80;
		memory[16'h7b54] <= 8'hc;
		memory[16'h7b55] <= 8'ha8;
		memory[16'h7b56] <= 8'h30;
		memory[16'h7b57] <= 8'h27;
		memory[16'h7b58] <= 8'h29;
		memory[16'h7b59] <= 8'h1a;
		memory[16'h7b5a] <= 8'h2b;
		memory[16'h7b5b] <= 8'h1b;
		memory[16'h7b5c] <= 8'h19;
		memory[16'h7b5d] <= 8'hd5;
		memory[16'h7b5e] <= 8'h83;
		memory[16'h7b5f] <= 8'h78;
		memory[16'h7b60] <= 8'hff;
		memory[16'h7b61] <= 8'h67;
		memory[16'h7b62] <= 8'hbd;
		memory[16'h7b63] <= 8'ha2;
		memory[16'h7b64] <= 8'hf9;
		memory[16'h7b65] <= 8'h1e;
		memory[16'h7b66] <= 8'hf0;
		memory[16'h7b67] <= 8'h4e;
		memory[16'h7b68] <= 8'h5f;
		memory[16'h7b69] <= 8'h24;
		memory[16'h7b6a] <= 8'hbf;
		memory[16'h7b6b] <= 8'he5;
		memory[16'h7b6c] <= 8'h6c;
		memory[16'h7b6d] <= 8'h64;
		memory[16'h7b6e] <= 8'h63;
		memory[16'h7b6f] <= 8'hda;
		memory[16'h7b70] <= 8'h27;
		memory[16'h7b71] <= 8'hee;
		memory[16'h7b72] <= 8'h5b;
		memory[16'h7b73] <= 8'h34;
		memory[16'h7b74] <= 8'h96;
		memory[16'h7b75] <= 8'h8b;
		memory[16'h7b76] <= 8'h5b;
		memory[16'h7b77] <= 8'hc0;
		memory[16'h7b78] <= 8'ha5;
		memory[16'h7b79] <= 8'h86;
		memory[16'h7b7a] <= 8'hdb;
		memory[16'h7b7b] <= 8'hbe;
		memory[16'h7b7c] <= 8'h5b;
		memory[16'h7b7d] <= 8'h5e;
		memory[16'h7b7e] <= 8'h36;
		memory[16'h7b7f] <= 8'h5a;
		memory[16'h7b80] <= 8'hc5;
		memory[16'h7b81] <= 8'hf4;
		memory[16'h7b82] <= 8'hfc;
		memory[16'h7b83] <= 8'hbe;
		memory[16'h7b84] <= 8'h12;
		memory[16'h7b85] <= 8'hec;
		memory[16'h7b86] <= 8'hd;
		memory[16'h7b87] <= 8'h71;
		memory[16'h7b88] <= 8'h11;
		memory[16'h7b89] <= 8'hcc;
		memory[16'h7b8a] <= 8'h56;
		memory[16'h7b8b] <= 8'h7d;
		memory[16'h7b8c] <= 8'h31;
		memory[16'h7b8d] <= 8'hba;
		memory[16'h7b8e] <= 8'h58;
		memory[16'h7b8f] <= 8'h58;
		memory[16'h7b90] <= 8'ha8;
		memory[16'h7b91] <= 8'hb3;
		memory[16'h7b92] <= 8'h8c;
		memory[16'h7b93] <= 8'h3f;
		memory[16'h7b94] <= 8'h3e;
		memory[16'h7b95] <= 8'he7;
		memory[16'h7b96] <= 8'hff;
		memory[16'h7b97] <= 8'he4;
		memory[16'h7b98] <= 8'h6d;
		memory[16'h7b99] <= 8'hda;
		memory[16'h7b9a] <= 8'ha2;
		memory[16'h7b9b] <= 8'hc9;
		memory[16'h7b9c] <= 8'h39;
		memory[16'h7b9d] <= 8'hd9;
		memory[16'h7b9e] <= 8'h23;
		memory[16'h7b9f] <= 8'hfe;
		memory[16'h7ba0] <= 8'hcd;
		memory[16'h7ba1] <= 8'h20;
		memory[16'h7ba2] <= 8'hbd;
		memory[16'h7ba3] <= 8'hdf;
		memory[16'h7ba4] <= 8'hc;
		memory[16'h7ba5] <= 8'hca;
		memory[16'h7ba6] <= 8'h51;
		memory[16'h7ba7] <= 8'h1d;
		memory[16'h7ba8] <= 8'h96;
		memory[16'h7ba9] <= 8'ha7;
		memory[16'h7baa] <= 8'h9b;
		memory[16'h7bab] <= 8'hc7;
		memory[16'h7bac] <= 8'h61;
		memory[16'h7bad] <= 8'hf3;
		memory[16'h7bae] <= 8'h20;
		memory[16'h7baf] <= 8'ha;
		memory[16'h7bb0] <= 8'ha6;
		memory[16'h7bb1] <= 8'hac;
		memory[16'h7bb2] <= 8'h49;
		memory[16'h7bb3] <= 8'he4;
		memory[16'h7bb4] <= 8'h94;
		memory[16'h7bb5] <= 8'h48;
		memory[16'h7bb6] <= 8'hc8;
		memory[16'h7bb7] <= 8'h1;
		memory[16'h7bb8] <= 8'h22;
		memory[16'h7bb9] <= 8'h6b;
		memory[16'h7bba] <= 8'hca;
		memory[16'h7bbb] <= 8'h5b;
		memory[16'h7bbc] <= 8'h44;
		memory[16'h7bbd] <= 8'hee;
		memory[16'h7bbe] <= 8'h5a;
		memory[16'h7bbf] <= 8'h11;
		memory[16'h7bc0] <= 8'he;
		memory[16'h7bc1] <= 8'h17;
		memory[16'h7bc2] <= 8'hf0;
		memory[16'h7bc3] <= 8'h1a;
		memory[16'h7bc4] <= 8'he1;
		memory[16'h7bc5] <= 8'h41;
		memory[16'h7bc6] <= 8'h38;
		memory[16'h7bc7] <= 8'h77;
		memory[16'h7bc8] <= 8'he9;
		memory[16'h7bc9] <= 8'hd3;
		memory[16'h7bca] <= 8'h3f;
		memory[16'h7bcb] <= 8'h4a;
		memory[16'h7bcc] <= 8'hc6;
		memory[16'h7bcd] <= 8'h5f;
		memory[16'h7bce] <= 8'h54;
		memory[16'h7bcf] <= 8'h6c;
		memory[16'h7bd0] <= 8'hb;
		memory[16'h7bd1] <= 8'h9d;
		memory[16'h7bd2] <= 8'h50;
		memory[16'h7bd3] <= 8'h9f;
		memory[16'h7bd4] <= 8'he5;
		memory[16'h7bd5] <= 8'h19;
		memory[16'h7bd6] <= 8'ha1;
		memory[16'h7bd7] <= 8'h8;
		memory[16'h7bd8] <= 8'h84;
		memory[16'h7bd9] <= 8'h6b;
		memory[16'h7bda] <= 8'h63;
		memory[16'h7bdb] <= 8'hc8;
		memory[16'h7bdc] <= 8'h59;
		memory[16'h7bdd] <= 8'hbd;
		memory[16'h7bde] <= 8'hd9;
		memory[16'h7bdf] <= 8'h67;
		memory[16'h7be0] <= 8'hd4;
		memory[16'h7be1] <= 8'hc9;
		memory[16'h7be2] <= 8'h82;
		memory[16'h7be3] <= 8'hb5;
		memory[16'h7be4] <= 8'hb;
		memory[16'h7be5] <= 8'hba;
		memory[16'h7be6] <= 8'h2d;
		memory[16'h7be7] <= 8'hf4;
		memory[16'h7be8] <= 8'h8d;
		memory[16'h7be9] <= 8'h6c;
		memory[16'h7bea] <= 8'h3e;
		memory[16'h7beb] <= 8'h53;
		memory[16'h7bec] <= 8'hcb;
		memory[16'h7bed] <= 8'h93;
		memory[16'h7bee] <= 8'hbf;
		memory[16'h7bef] <= 8'hd6;
		memory[16'h7bf0] <= 8'h30;
		memory[16'h7bf1] <= 8'hf;
		memory[16'h7bf2] <= 8'h76;
		memory[16'h7bf3] <= 8'h16;
		memory[16'h7bf4] <= 8'h28;
		memory[16'h7bf5] <= 8'h17;
		memory[16'h7bf6] <= 8'h1e;
		memory[16'h7bf7] <= 8'hac;
		memory[16'h7bf8] <= 8'h82;
		memory[16'h7bf9] <= 8'h81;
		memory[16'h7bfa] <= 8'h74;
		memory[16'h7bfb] <= 8'hdc;
		memory[16'h7bfc] <= 8'h3f;
		memory[16'h7bfd] <= 8'h4d;
		memory[16'h7bfe] <= 8'h43;
		memory[16'h7bff] <= 8'h13;
		memory[16'h7c00] <= 8'h17;
		memory[16'h7c01] <= 8'hc5;
		memory[16'h7c02] <= 8'hc9;
		memory[16'h7c03] <= 8'h22;
		memory[16'h7c04] <= 8'h7f;
		memory[16'h7c05] <= 8'hf6;
		memory[16'h7c06] <= 8'h16;
		memory[16'h7c07] <= 8'hc;
		memory[16'h7c08] <= 8'h62;
		memory[16'h7c09] <= 8'h54;
		memory[16'h7c0a] <= 8'h5f;
		memory[16'h7c0b] <= 8'h2d;
		memory[16'h7c0c] <= 8'he7;
		memory[16'h7c0d] <= 8'h1e;
		memory[16'h7c0e] <= 8'h3;
		memory[16'h7c0f] <= 8'h18;
		memory[16'h7c10] <= 8'h2e;
		memory[16'h7c11] <= 8'h79;
		memory[16'h7c12] <= 8'h2e;
		memory[16'h7c13] <= 8'h56;
		memory[16'h7c14] <= 8'h90;
		memory[16'h7c15] <= 8'h4c;
		memory[16'h7c16] <= 8'h3;
		memory[16'h7c17] <= 8'h13;
		memory[16'h7c18] <= 8'hcd;
		memory[16'h7c19] <= 8'h77;
		memory[16'h7c1a] <= 8'hef;
		memory[16'h7c1b] <= 8'hc;
		memory[16'h7c1c] <= 8'hc5;
		memory[16'h7c1d] <= 8'h32;
		memory[16'h7c1e] <= 8'h20;
		memory[16'h7c1f] <= 8'hdc;
		memory[16'h7c20] <= 8'hf8;
		memory[16'h7c21] <= 8'he9;
		memory[16'h7c22] <= 8'hfe;
		memory[16'h7c23] <= 8'h77;
		memory[16'h7c24] <= 8'hdf;
		memory[16'h7c25] <= 8'h14;
		memory[16'h7c26] <= 8'h84;
		memory[16'h7c27] <= 8'h41;
		memory[16'h7c28] <= 8'h68;
		memory[16'h7c29] <= 8'he3;
		memory[16'h7c2a] <= 8'h6e;
		memory[16'h7c2b] <= 8'h50;
		memory[16'h7c2c] <= 8'h2;
		memory[16'h7c2d] <= 8'h71;
		memory[16'h7c2e] <= 8'h68;
		memory[16'h7c2f] <= 8'h30;
		memory[16'h7c30] <= 8'heb;
		memory[16'h7c31] <= 8'h96;
		memory[16'h7c32] <= 8'h86;
		memory[16'h7c33] <= 8'h7b;
		memory[16'h7c34] <= 8'he2;
		memory[16'h7c35] <= 8'h89;
		memory[16'h7c36] <= 8'h8e;
		memory[16'h7c37] <= 8'haf;
		memory[16'h7c38] <= 8'h1;
		memory[16'h7c39] <= 8'h7d;
		memory[16'h7c3a] <= 8'hbc;
		memory[16'h7c3b] <= 8'hc6;
		memory[16'h7c3c] <= 8'hb0;
		memory[16'h7c3d] <= 8'hdc;
		memory[16'h7c3e] <= 8'ha2;
		memory[16'h7c3f] <= 8'ha8;
		memory[16'h7c40] <= 8'hc5;
		memory[16'h7c41] <= 8'ha0;
		memory[16'h7c42] <= 8'h1f;
		memory[16'h7c43] <= 8'ha4;
		memory[16'h7c44] <= 8'hb4;
		memory[16'h7c45] <= 8'ha3;
		memory[16'h7c46] <= 8'he5;
		memory[16'h7c47] <= 8'h1c;
		memory[16'h7c48] <= 8'h87;
		memory[16'h7c49] <= 8'h53;
		memory[16'h7c4a] <= 8'h6c;
		memory[16'h7c4b] <= 8'h89;
		memory[16'h7c4c] <= 8'hc4;
		memory[16'h7c4d] <= 8'hd4;
		memory[16'h7c4e] <= 8'hb9;
		memory[16'h7c4f] <= 8'haf;
		memory[16'h7c50] <= 8'h6a;
		memory[16'h7c51] <= 8'h3f;
		memory[16'h7c52] <= 8'h2b;
		memory[16'h7c53] <= 8'h4c;
		memory[16'h7c54] <= 8'hc9;
		memory[16'h7c55] <= 8'hb9;
		memory[16'h7c56] <= 8'hfc;
		memory[16'h7c57] <= 8'hca;
		memory[16'h7c58] <= 8'h37;
		memory[16'h7c59] <= 8'hb8;
		memory[16'h7c5a] <= 8'h90;
		memory[16'h7c5b] <= 8'he7;
		memory[16'h7c5c] <= 8'h94;
		memory[16'h7c5d] <= 8'h32;
		memory[16'h7c5e] <= 8'h8f;
		memory[16'h7c5f] <= 8'h59;
		memory[16'h7c60] <= 8'hd2;
		memory[16'h7c61] <= 8'hae;
		memory[16'h7c62] <= 8'hfd;
		memory[16'h7c63] <= 8'h86;
		memory[16'h7c64] <= 8'h52;
		memory[16'h7c65] <= 8'he2;
		memory[16'h7c66] <= 8'ha2;
		memory[16'h7c67] <= 8'hd9;
		memory[16'h7c68] <= 8'h35;
		memory[16'h7c69] <= 8'hf;
		memory[16'h7c6a] <= 8'h62;
		memory[16'h7c6b] <= 8'hf9;
		memory[16'h7c6c] <= 8'he3;
		memory[16'h7c6d] <= 8'h1b;
		memory[16'h7c6e] <= 8'ha9;
		memory[16'h7c6f] <= 8'h4e;
		memory[16'h7c70] <= 8'h5a;
		memory[16'h7c71] <= 8'hd4;
		memory[16'h7c72] <= 8'h9a;
		memory[16'h7c73] <= 8'h23;
		memory[16'h7c74] <= 8'h8d;
		memory[16'h7c75] <= 8'h96;
		memory[16'h7c76] <= 8'hed;
		memory[16'h7c77] <= 8'hc4;
		memory[16'h7c78] <= 8'h4e;
		memory[16'h7c79] <= 8'h7d;
		memory[16'h7c7a] <= 8'hab;
		memory[16'h7c7b] <= 8'he2;
		memory[16'h7c7c] <= 8'haf;
		memory[16'h7c7d] <= 8'h3a;
		memory[16'h7c7e] <= 8'h3b;
		memory[16'h7c7f] <= 8'h81;
		memory[16'h7c80] <= 8'he9;
		memory[16'h7c81] <= 8'h38;
		memory[16'h7c82] <= 8'h7;
		memory[16'h7c83] <= 8'h3b;
		memory[16'h7c84] <= 8'h1a;
		memory[16'h7c85] <= 8'haa;
		memory[16'h7c86] <= 8'h14;
		memory[16'h7c87] <= 8'h4f;
		memory[16'h7c88] <= 8'hb9;
		memory[16'h7c89] <= 8'h76;
		memory[16'h7c8a] <= 8'h49;
		memory[16'h7c8b] <= 8'h9c;
		memory[16'h7c8c] <= 8'h91;
		memory[16'h7c8d] <= 8'hf2;
		memory[16'h7c8e] <= 8'hea;
		memory[16'h7c8f] <= 8'heb;
		memory[16'h7c90] <= 8'hc6;
		memory[16'h7c91] <= 8'h85;
		memory[16'h7c92] <= 8'hf;
		memory[16'h7c93] <= 8'h53;
		memory[16'h7c94] <= 8'h1b;
		memory[16'h7c95] <= 8'hfc;
		memory[16'h7c96] <= 8'h18;
		memory[16'h7c97] <= 8'h6a;
		memory[16'h7c98] <= 8'h7a;
		memory[16'h7c99] <= 8'hc3;
		memory[16'h7c9a] <= 8'h4c;
		memory[16'h7c9b] <= 8'h29;
		memory[16'h7c9c] <= 8'hfe;
		memory[16'h7c9d] <= 8'h88;
		memory[16'h7c9e] <= 8'hab;
		memory[16'h7c9f] <= 8'he7;
		memory[16'h7ca0] <= 8'hc0;
		memory[16'h7ca1] <= 8'hb2;
		memory[16'h7ca2] <= 8'h22;
		memory[16'h7ca3] <= 8'hdb;
		memory[16'h7ca4] <= 8'h5c;
		memory[16'h7ca5] <= 8'h36;
		memory[16'h7ca6] <= 8'h2a;
		memory[16'h7ca7] <= 8'h15;
		memory[16'h7ca8] <= 8'hac;
		memory[16'h7ca9] <= 8'h73;
		memory[16'h7caa] <= 8'hb2;
		memory[16'h7cab] <= 8'h3d;
		memory[16'h7cac] <= 8'h65;
		memory[16'h7cad] <= 8'h9c;
		memory[16'h7cae] <= 8'h28;
		memory[16'h7caf] <= 8'h2b;
		memory[16'h7cb0] <= 8'h21;
		memory[16'h7cb1] <= 8'h37;
		memory[16'h7cb2] <= 8'h7f;
		memory[16'h7cb3] <= 8'h3d;
		memory[16'h7cb4] <= 8'h34;
		memory[16'h7cb5] <= 8'h97;
		memory[16'h7cb6] <= 8'ha7;
		memory[16'h7cb7] <= 8'hae;
		memory[16'h7cb8] <= 8'h5a;
		memory[16'h7cb9] <= 8'hf3;
		memory[16'h7cba] <= 8'hd7;
		memory[16'h7cbb] <= 8'h58;
		memory[16'h7cbc] <= 8'h7b;
		memory[16'h7cbd] <= 8'h82;
		memory[16'h7cbe] <= 8'h3f;
		memory[16'h7cbf] <= 8'h3c;
		memory[16'h7cc0] <= 8'h35;
		memory[16'h7cc1] <= 8'h61;
		memory[16'h7cc2] <= 8'h17;
		memory[16'h7cc3] <= 8'h91;
		memory[16'h7cc4] <= 8'h97;
		memory[16'h7cc5] <= 8'h41;
		memory[16'h7cc6] <= 8'ha7;
		memory[16'h7cc7] <= 8'h43;
		memory[16'h7cc8] <= 8'hb5;
		memory[16'h7cc9] <= 8'h59;
		memory[16'h7cca] <= 8'h80;
		memory[16'h7ccb] <= 8'h1a;
		memory[16'h7ccc] <= 8'hf5;
		memory[16'h7ccd] <= 8'ha9;
		memory[16'h7cce] <= 8'h46;
		memory[16'h7ccf] <= 8'h17;
		memory[16'h7cd0] <= 8'he0;
		memory[16'h7cd1] <= 8'hc5;
		memory[16'h7cd2] <= 8'h54;
		memory[16'h7cd3] <= 8'h14;
		memory[16'h7cd4] <= 8'h5c;
		memory[16'h7cd5] <= 8'hfb;
		memory[16'h7cd6] <= 8'hc2;
		memory[16'h7cd7] <= 8'hb6;
		memory[16'h7cd8] <= 8'hee;
		memory[16'h7cd9] <= 8'h9a;
		memory[16'h7cda] <= 8'hf;
		memory[16'h7cdb] <= 8'h6a;
		memory[16'h7cdc] <= 8'h1c;
		memory[16'h7cdd] <= 8'h4e;
		memory[16'h7cde] <= 8'ha6;
		memory[16'h7cdf] <= 8'h51;
		memory[16'h7ce0] <= 8'hb0;
		memory[16'h7ce1] <= 8'hbd;
		memory[16'h7ce2] <= 8'he3;
		memory[16'h7ce3] <= 8'h47;
		memory[16'h7ce4] <= 8'hfe;
		memory[16'h7ce5] <= 8'h8a;
		memory[16'h7ce6] <= 8'h8b;
		memory[16'h7ce7] <= 8'hb3;
		memory[16'h7ce8] <= 8'he3;
		memory[16'h7ce9] <= 8'hb;
		memory[16'h7cea] <= 8'hce;
		memory[16'h7ceb] <= 8'hd8;
		memory[16'h7cec] <= 8'hb4;
		memory[16'h7ced] <= 8'h14;
		memory[16'h7cee] <= 8'hef;
		memory[16'h7cef] <= 8'h95;
		memory[16'h7cf0] <= 8'hd9;
		memory[16'h7cf1] <= 8'h43;
		memory[16'h7cf2] <= 8'ha9;
		memory[16'h7cf3] <= 8'h35;
		memory[16'h7cf4] <= 8'h3e;
		memory[16'h7cf5] <= 8'h6c;
		memory[16'h7cf6] <= 8'heb;
		memory[16'h7cf7] <= 8'h2d;
		memory[16'h7cf8] <= 8'h6;
		memory[16'h7cf9] <= 8'hfa;
		memory[16'h7cfa] <= 8'h97;
		memory[16'h7cfb] <= 8'h22;
		memory[16'h7cfc] <= 8'h49;
		memory[16'h7cfd] <= 8'h3d;
		memory[16'h7cfe] <= 8'h74;
		memory[16'h7cff] <= 8'hf9;
		memory[16'h7d00] <= 8'hfa;
		memory[16'h7d01] <= 8'h57;
		memory[16'h7d02] <= 8'h40;
		memory[16'h7d03] <= 8'hf8;
		memory[16'h7d04] <= 8'he1;
		memory[16'h7d05] <= 8'hcb;
		memory[16'h7d06] <= 8'hac;
		memory[16'h7d07] <= 8'hc4;
		memory[16'h7d08] <= 8'hd7;
		memory[16'h7d09] <= 8'h7a;
		memory[16'h7d0a] <= 8'h9c;
		memory[16'h7d0b] <= 8'h8b;
		memory[16'h7d0c] <= 8'h8e;
		memory[16'h7d0d] <= 8'h8c;
		memory[16'h7d0e] <= 8'h20;
		memory[16'h7d0f] <= 8'h67;
		memory[16'h7d10] <= 8'hcf;
		memory[16'h7d11] <= 8'hca;
		memory[16'h7d12] <= 8'h9c;
		memory[16'h7d13] <= 8'he;
		memory[16'h7d14] <= 8'h36;
		memory[16'h7d15] <= 8'h87;
		memory[16'h7d16] <= 8'h3b;
		memory[16'h7d17] <= 8'h3c;
		memory[16'h7d18] <= 8'h82;
		memory[16'h7d19] <= 8'hd2;
		memory[16'h7d1a] <= 8'h5e;
		memory[16'h7d1b] <= 8'hcb;
		memory[16'h7d1c] <= 8'hf;
		memory[16'h7d1d] <= 8'hd2;
		memory[16'h7d1e] <= 8'hc4;
		memory[16'h7d1f] <= 8'h9;
		memory[16'h7d20] <= 8'h29;
		memory[16'h7d21] <= 8'h4;
		memory[16'h7d22] <= 8'h1;
		memory[16'h7d23] <= 8'ha;
		memory[16'h7d24] <= 8'hd0;
		memory[16'h7d25] <= 8'had;
		memory[16'h7d26] <= 8'hce;
		memory[16'h7d27] <= 8'ha7;
		memory[16'h7d28] <= 8'h27;
		memory[16'h7d29] <= 8'h6b;
		memory[16'h7d2a] <= 8'h32;
		memory[16'h7d2b] <= 8'hb5;
		memory[16'h7d2c] <= 8'hf7;
		memory[16'h7d2d] <= 8'h53;
		memory[16'h7d2e] <= 8'h1c;
		memory[16'h7d2f] <= 8'hc6;
		memory[16'h7d30] <= 8'h1d;
		memory[16'h7d31] <= 8'hb8;
		memory[16'h7d32] <= 8'hd4;
		memory[16'h7d33] <= 8'h53;
		memory[16'h7d34] <= 8'h40;
		memory[16'h7d35] <= 8'hf;
		memory[16'h7d36] <= 8'h8f;
		memory[16'h7d37] <= 8'hc2;
		memory[16'h7d38] <= 8'he1;
		memory[16'h7d39] <= 8'hed;
		memory[16'h7d3a] <= 8'h8d;
		memory[16'h7d3b] <= 8'hf0;
		memory[16'h7d3c] <= 8'hc0;
		memory[16'h7d3d] <= 8'h51;
		memory[16'h7d3e] <= 8'hf9;
		memory[16'h7d3f] <= 8'he9;
		memory[16'h7d40] <= 8'h55;
		memory[16'h7d41] <= 8'hfb;
		memory[16'h7d42] <= 8'hf4;
		memory[16'h7d43] <= 8'h25;
		memory[16'h7d44] <= 8'ha8;
		memory[16'h7d45] <= 8'hc2;
		memory[16'h7d46] <= 8'hcc;
		memory[16'h7d47] <= 8'hd0;
		memory[16'h7d48] <= 8'h2d;
		memory[16'h7d49] <= 8'hff;
		memory[16'h7d4a] <= 8'h85;
		memory[16'h7d4b] <= 8'h24;
		memory[16'h7d4c] <= 8'h52;
		memory[16'h7d4d] <= 8'ha2;
		memory[16'h7d4e] <= 8'heb;
		memory[16'h7d4f] <= 8'h6f;
		memory[16'h7d50] <= 8'h5a;
		memory[16'h7d51] <= 8'hbf;
		memory[16'h7d52] <= 8'hc2;
		memory[16'h7d53] <= 8'h9a;
		memory[16'h7d54] <= 8'hcf;
		memory[16'h7d55] <= 8'h51;
		memory[16'h7d56] <= 8'h5c;
		memory[16'h7d57] <= 8'hb0;
		memory[16'h7d58] <= 8'h3e;
		memory[16'h7d59] <= 8'he9;
		memory[16'h7d5a] <= 8'ha1;
		memory[16'h7d5b] <= 8'hfe;
		memory[16'h7d5c] <= 8'h3a;
		memory[16'h7d5d] <= 8'h9a;
		memory[16'h7d5e] <= 8'he8;
		memory[16'h7d5f] <= 8'h90;
		memory[16'h7d60] <= 8'h95;
		memory[16'h7d61] <= 8'hdc;
		memory[16'h7d62] <= 8'hb5;
		memory[16'h7d63] <= 8'h3e;
		memory[16'h7d64] <= 8'h9e;
		memory[16'h7d65] <= 8'h82;
		memory[16'h7d66] <= 8'he;
		memory[16'h7d67] <= 8'hcc;
		memory[16'h7d68] <= 8'h81;
		memory[16'h7d69] <= 8'h93;
		memory[16'h7d6a] <= 8'hf0;
		memory[16'h7d6b] <= 8'hd3;
		memory[16'h7d6c] <= 8'h35;
		memory[16'h7d6d] <= 8'hdb;
		memory[16'h7d6e] <= 8'h42;
		memory[16'h7d6f] <= 8'h90;
		memory[16'h7d70] <= 8'h9b;
		memory[16'h7d71] <= 8'h4;
		memory[16'h7d72] <= 8'h2a;
		memory[16'h7d73] <= 8'h6a;
		memory[16'h7d74] <= 8'h55;
		memory[16'h7d75] <= 8'h87;
		memory[16'h7d76] <= 8'h1a;
		memory[16'h7d77] <= 8'h93;
		memory[16'h7d78] <= 8'h70;
		memory[16'h7d79] <= 8'hbb;
		memory[16'h7d7a] <= 8'h92;
		memory[16'h7d7b] <= 8'hab;
		memory[16'h7d7c] <= 8'h56;
		memory[16'h7d7d] <= 8'h7a;
		memory[16'h7d7e] <= 8'h3b;
		memory[16'h7d7f] <= 8'heb;
		memory[16'h7d80] <= 8'h56;
		memory[16'h7d81] <= 8'hf0;
		memory[16'h7d82] <= 8'h29;
		memory[16'h7d83] <= 8'hf4;
		memory[16'h7d84] <= 8'h72;
		memory[16'h7d85] <= 8'h37;
		memory[16'h7d86] <= 8'hc0;
		memory[16'h7d87] <= 8'hf3;
		memory[16'h7d88] <= 8'hcb;
		memory[16'h7d89] <= 8'hb1;
		memory[16'h7d8a] <= 8'hc6;
		memory[16'h7d8b] <= 8'h0;
		memory[16'h7d8c] <= 8'h8c;
		memory[16'h7d8d] <= 8'h8;
		memory[16'h7d8e] <= 8'h90;
		memory[16'h7d8f] <= 8'h27;
		memory[16'h7d90] <= 8'hc;
		memory[16'h7d91] <= 8'hbb;
		memory[16'h7d92] <= 8'h91;
		memory[16'h7d93] <= 8'h61;
		memory[16'h7d94] <= 8'h42;
		memory[16'h7d95] <= 8'hac;
		memory[16'h7d96] <= 8'hf5;
		memory[16'h7d97] <= 8'hb2;
		memory[16'h7d98] <= 8'h67;
		memory[16'h7d99] <= 8'h87;
		memory[16'h7d9a] <= 8'h5d;
		memory[16'h7d9b] <= 8'hbd;
		memory[16'h7d9c] <= 8'h1;
		memory[16'h7d9d] <= 8'h98;
		memory[16'h7d9e] <= 8'ha9;
		memory[16'h7d9f] <= 8'h57;
		memory[16'h7da0] <= 8'h89;
		memory[16'h7da1] <= 8'hd2;
		memory[16'h7da2] <= 8'h4b;
		memory[16'h7da3] <= 8'hfb;
		memory[16'h7da4] <= 8'ha;
		memory[16'h7da5] <= 8'hc;
		memory[16'h7da6] <= 8'hef;
		memory[16'h7da7] <= 8'hd5;
		memory[16'h7da8] <= 8'hbd;
		memory[16'h7da9] <= 8'hb5;
		memory[16'h7daa] <= 8'hd5;
		memory[16'h7dab] <= 8'h49;
		memory[16'h7dac] <= 8'hbe;
		memory[16'h7dad] <= 8'h66;
		memory[16'h7dae] <= 8'h71;
		memory[16'h7daf] <= 8'hca;
		memory[16'h7db0] <= 8'h21;
		memory[16'h7db1] <= 8'h2;
		memory[16'h7db2] <= 8'h2c;
		memory[16'h7db3] <= 8'h63;
		memory[16'h7db4] <= 8'hae;
		memory[16'h7db5] <= 8'h21;
		memory[16'h7db6] <= 8'h15;
		memory[16'h7db7] <= 8'h16;
		memory[16'h7db8] <= 8'ha8;
		memory[16'h7db9] <= 8'h73;
		memory[16'h7dba] <= 8'hd3;
		memory[16'h7dbb] <= 8'ha9;
		memory[16'h7dbc] <= 8'hb;
		memory[16'h7dbd] <= 8'h7c;
		memory[16'h7dbe] <= 8'h0;
		memory[16'h7dbf] <= 8'h94;
		memory[16'h7dc0] <= 8'h4f;
		memory[16'h7dc1] <= 8'h4b;
		memory[16'h7dc2] <= 8'h90;
		memory[16'h7dc3] <= 8'h59;
		memory[16'h7dc4] <= 8'h57;
		memory[16'h7dc5] <= 8'h7f;
		memory[16'h7dc6] <= 8'h2e;
		memory[16'h7dc7] <= 8'h14;
		memory[16'h7dc8] <= 8'h34;
		memory[16'h7dc9] <= 8'h3;
		memory[16'h7dca] <= 8'h5e;
		memory[16'h7dcb] <= 8'hf2;
		memory[16'h7dcc] <= 8'h69;
		memory[16'h7dcd] <= 8'hcf;
		memory[16'h7dce] <= 8'hbd;
		memory[16'h7dcf] <= 8'h8a;
		memory[16'h7dd0] <= 8'hd1;
		memory[16'h7dd1] <= 8'he9;
		memory[16'h7dd2] <= 8'hed;
		memory[16'h7dd3] <= 8'h80;
		memory[16'h7dd4] <= 8'ha;
		memory[16'h7dd5] <= 8'h3;
		memory[16'h7dd6] <= 8'h96;
		memory[16'h7dd7] <= 8'hb2;
		memory[16'h7dd8] <= 8'h76;
		memory[16'h7dd9] <= 8'h69;
		memory[16'h7dda] <= 8'h5b;
		memory[16'h7ddb] <= 8'h81;
		memory[16'h7ddc] <= 8'he6;
		memory[16'h7ddd] <= 8'h5b;
		memory[16'h7dde] <= 8'h16;
		memory[16'h7ddf] <= 8'h35;
		memory[16'h7de0] <= 8'ha6;
		memory[16'h7de1] <= 8'ha6;
		memory[16'h7de2] <= 8'h8e;
		memory[16'h7de3] <= 8'hfe;
		memory[16'h7de4] <= 8'h25;
		memory[16'h7de5] <= 8'hbc;
		memory[16'h7de6] <= 8'h12;
		memory[16'h7de7] <= 8'h59;
		memory[16'h7de8] <= 8'hbf;
		memory[16'h7de9] <= 8'h70;
		memory[16'h7dea] <= 8'h4c;
		memory[16'h7deb] <= 8'h29;
		memory[16'h7dec] <= 8'h3f;
		memory[16'h7ded] <= 8'h9;
		memory[16'h7dee] <= 8'hb3;
		memory[16'h7def] <= 8'h11;
		memory[16'h7df0] <= 8'hf2;
		memory[16'h7df1] <= 8'ha1;
		memory[16'h7df2] <= 8'h91;
		memory[16'h7df3] <= 8'hfc;
		memory[16'h7df4] <= 8'ha4;
		memory[16'h7df5] <= 8'h27;
		memory[16'h7df6] <= 8'hae;
		memory[16'h7df7] <= 8'h1a;
		memory[16'h7df8] <= 8'h90;
		memory[16'h7df9] <= 8'h9;
		memory[16'h7dfa] <= 8'h9b;
		memory[16'h7dfb] <= 8'h76;
		memory[16'h7dfc] <= 8'h64;
		memory[16'h7dfd] <= 8'hb1;
		memory[16'h7dfe] <= 8'hab;
		memory[16'h7dff] <= 8'ha;
		memory[16'h7e00] <= 8'h57;
		memory[16'h7e01] <= 8'h39;
		memory[16'h7e02] <= 8'h8;
		memory[16'h7e03] <= 8'h7c;
		memory[16'h7e04] <= 8'hf5;
		memory[16'h7e05] <= 8'h1b;
		memory[16'h7e06] <= 8'hd6;
		memory[16'h7e07] <= 8'hb5;
		memory[16'h7e08] <= 8'h8b;
		memory[16'h7e09] <= 8'h22;
		memory[16'h7e0a] <= 8'hde;
		memory[16'h7e0b] <= 8'hcb;
		memory[16'h7e0c] <= 8'h2b;
		memory[16'h7e0d] <= 8'h91;
		memory[16'h7e0e] <= 8'hdc;
		memory[16'h7e0f] <= 8'h1d;
		memory[16'h7e10] <= 8'h32;
		memory[16'h7e11] <= 8'h6d;
		memory[16'h7e12] <= 8'h19;
		memory[16'h7e13] <= 8'hd6;
		memory[16'h7e14] <= 8'h94;
		memory[16'h7e15] <= 8'hc7;
		memory[16'h7e16] <= 8'hf0;
		memory[16'h7e17] <= 8'h24;
		memory[16'h7e18] <= 8'hd0;
		memory[16'h7e19] <= 8'h8c;
		memory[16'h7e1a] <= 8'h9b;
		memory[16'h7e1b] <= 8'h34;
		memory[16'h7e1c] <= 8'h3d;
		memory[16'h7e1d] <= 8'h46;
		memory[16'h7e1e] <= 8'h3e;
		memory[16'h7e1f] <= 8'h95;
		memory[16'h7e20] <= 8'h80;
		memory[16'h7e21] <= 8'h47;
		memory[16'h7e22] <= 8'h11;
		memory[16'h7e23] <= 8'h75;
		memory[16'h7e24] <= 8'h62;
		memory[16'h7e25] <= 8'he7;
		memory[16'h7e26] <= 8'h2a;
		memory[16'h7e27] <= 8'hed;
		memory[16'h7e28] <= 8'h9;
		memory[16'h7e29] <= 8'h8;
		memory[16'h7e2a] <= 8'hb8;
		memory[16'h7e2b] <= 8'h34;
		memory[16'h7e2c] <= 8'h9a;
		memory[16'h7e2d] <= 8'h94;
		memory[16'h7e2e] <= 8'h51;
		memory[16'h7e2f] <= 8'hcc;
		memory[16'h7e30] <= 8'h1;
		memory[16'h7e31] <= 8'h6a;
		memory[16'h7e32] <= 8'ha3;
		memory[16'h7e33] <= 8'h95;
		memory[16'h7e34] <= 8'h31;
		memory[16'h7e35] <= 8'h93;
		memory[16'h7e36] <= 8'hba;
		memory[16'h7e37] <= 8'h1;
		memory[16'h7e38] <= 8'h1f;
		memory[16'h7e39] <= 8'h55;
		memory[16'h7e3a] <= 8'h35;
		memory[16'h7e3b] <= 8'h5d;
		memory[16'h7e3c] <= 8'h9b;
		memory[16'h7e3d] <= 8'h74;
		memory[16'h7e3e] <= 8'hf2;
		memory[16'h7e3f] <= 8'h1b;
		memory[16'h7e40] <= 8'hbb;
		memory[16'h7e41] <= 8'h3;
		memory[16'h7e42] <= 8'h91;
		memory[16'h7e43] <= 8'h1d;
		memory[16'h7e44] <= 8'heb;
		memory[16'h7e45] <= 8'hbb;
		memory[16'h7e46] <= 8'ha;
		memory[16'h7e47] <= 8'hf4;
		memory[16'h7e48] <= 8'hc4;
		memory[16'h7e49] <= 8'hc3;
		memory[16'h7e4a] <= 8'h29;
		memory[16'h7e4b] <= 8'h5e;
		memory[16'h7e4c] <= 8'h57;
		memory[16'h7e4d] <= 8'h7a;
		memory[16'h7e4e] <= 8'h2a;
		memory[16'h7e4f] <= 8'h59;
		memory[16'h7e50] <= 8'he5;
		memory[16'h7e51] <= 8'hcd;
		memory[16'h7e52] <= 8'hee;
		memory[16'h7e53] <= 8'h16;
		memory[16'h7e54] <= 8'h61;
		memory[16'h7e55] <= 8'ha8;
		memory[16'h7e56] <= 8'h18;
		memory[16'h7e57] <= 8'h80;
		memory[16'h7e58] <= 8'hfd;
		memory[16'h7e59] <= 8'h4d;
		memory[16'h7e5a] <= 8'hdd;
		memory[16'h7e5b] <= 8'h99;
		memory[16'h7e5c] <= 8'hc1;
		memory[16'h7e5d] <= 8'hcf;
		memory[16'h7e5e] <= 8'hb4;
		memory[16'h7e5f] <= 8'h7c;
		memory[16'h7e60] <= 8'hd3;
		memory[16'h7e61] <= 8'h45;
		memory[16'h7e62] <= 8'h99;
		memory[16'h7e63] <= 8'hbe;
		memory[16'h7e64] <= 8'h1;
		memory[16'h7e65] <= 8'ha4;
		memory[16'h7e66] <= 8'hb2;
		memory[16'h7e67] <= 8'hc5;
		memory[16'h7e68] <= 8'h67;
		memory[16'h7e69] <= 8'hdb;
		memory[16'h7e6a] <= 8'h23;
		memory[16'h7e6b] <= 8'hbe;
		memory[16'h7e6c] <= 8'h56;
		memory[16'h7e6d] <= 8'h4d;
		memory[16'h7e6e] <= 8'h17;
		memory[16'h7e6f] <= 8'h3b;
		memory[16'h7e70] <= 8'h1b;
		memory[16'h7e71] <= 8'h6;
		memory[16'h7e72] <= 8'h51;
		memory[16'h7e73] <= 8'h7c;
		memory[16'h7e74] <= 8'hae;
		memory[16'h7e75] <= 8'h69;
		memory[16'h7e76] <= 8'hfc;
		memory[16'h7e77] <= 8'hac;
		memory[16'h7e78] <= 8'hb7;
		memory[16'h7e79] <= 8'hda;
		memory[16'h7e7a] <= 8'h45;
		memory[16'h7e7b] <= 8'h78;
		memory[16'h7e7c] <= 8'ha9;
		memory[16'h7e7d] <= 8'hf9;
		memory[16'h7e7e] <= 8'hf5;
		memory[16'h7e7f] <= 8'h7c;
		memory[16'h7e80] <= 8'h3f;
		memory[16'h7e81] <= 8'h8e;
		memory[16'h7e82] <= 8'h3a;
		memory[16'h7e83] <= 8'h40;
		memory[16'h7e84] <= 8'h32;
		memory[16'h7e85] <= 8'hed;
		memory[16'h7e86] <= 8'h5;
		memory[16'h7e87] <= 8'h99;
		memory[16'h7e88] <= 8'hc8;
		memory[16'h7e89] <= 8'h28;
		memory[16'h7e8a] <= 8'h58;
		memory[16'h7e8b] <= 8'h1e;
		memory[16'h7e8c] <= 8'h75;
		memory[16'h7e8d] <= 8'h6f;
		memory[16'h7e8e] <= 8'h59;
		memory[16'h7e8f] <= 8'h90;
		memory[16'h7e90] <= 8'h75;
		memory[16'h7e91] <= 8'hab;
		memory[16'h7e92] <= 8'hc;
		memory[16'h7e93] <= 8'h24;
		memory[16'h7e94] <= 8'h14;
		memory[16'h7e95] <= 8'h9;
		memory[16'h7e96] <= 8'hd0;
		memory[16'h7e97] <= 8'hcb;
		memory[16'h7e98] <= 8'he3;
		memory[16'h7e99] <= 8'h15;
		memory[16'h7e9a] <= 8'h44;
		memory[16'h7e9b] <= 8'h8c;
		memory[16'h7e9c] <= 8'he;
		memory[16'h7e9d] <= 8'h39;
		memory[16'h7e9e] <= 8'h9;
		memory[16'h7e9f] <= 8'h4d;
		memory[16'h7ea0] <= 8'hc7;
		memory[16'h7ea1] <= 8'h43;
		memory[16'h7ea2] <= 8'h8d;
		memory[16'h7ea3] <= 8'hfa;
		memory[16'h7ea4] <= 8'h30;
		memory[16'h7ea5] <= 8'h92;
		memory[16'h7ea6] <= 8'h93;
		memory[16'h7ea7] <= 8'hf9;
		memory[16'h7ea8] <= 8'hba;
		memory[16'h7ea9] <= 8'heb;
		memory[16'h7eaa] <= 8'h17;
		memory[16'h7eab] <= 8'h30;
		memory[16'h7eac] <= 8'h5b;
		memory[16'h7ead] <= 8'h71;
		memory[16'h7eae] <= 8'hc0;
		memory[16'h7eaf] <= 8'hd0;
		memory[16'h7eb0] <= 8'h1c;
		memory[16'h7eb1] <= 8'hcd;
		memory[16'h7eb2] <= 8'hf4;
		memory[16'h7eb3] <= 8'h30;
		memory[16'h7eb4] <= 8'hd6;
		memory[16'h7eb5] <= 8'hc4;
		memory[16'h7eb6] <= 8'hfc;
		memory[16'h7eb7] <= 8'hb9;
		memory[16'h7eb8] <= 8'hd9;
		memory[16'h7eb9] <= 8'h40;
		memory[16'h7eba] <= 8'h45;
		memory[16'h7ebb] <= 8'he8;
		memory[16'h7ebc] <= 8'h79;
		memory[16'h7ebd] <= 8'h4e;
		memory[16'h7ebe] <= 8'h35;
		memory[16'h7ebf] <= 8'h40;
		memory[16'h7ec0] <= 8'h92;
		memory[16'h7ec1] <= 8'hc3;
		memory[16'h7ec2] <= 8'h3a;
		memory[16'h7ec3] <= 8'hc2;
		memory[16'h7ec4] <= 8'h55;
		memory[16'h7ec5] <= 8'hce;
		memory[16'h7ec6] <= 8'hbb;
		memory[16'h7ec7] <= 8'h10;
		memory[16'h7ec8] <= 8'hb9;
		memory[16'h7ec9] <= 8'hd3;
		memory[16'h7eca] <= 8'h40;
		memory[16'h7ecb] <= 8'h14;
		memory[16'h7ecc] <= 8'h44;
		memory[16'h7ecd] <= 8'h0;
		memory[16'h7ece] <= 8'he5;
		memory[16'h7ecf] <= 8'h60;
		memory[16'h7ed0] <= 8'hcd;
		memory[16'h7ed1] <= 8'hd9;
		memory[16'h7ed2] <= 8'h90;
		memory[16'h7ed3] <= 8'ha3;
		memory[16'h7ed4] <= 8'h9e;
		memory[16'h7ed5] <= 8'h8c;
		memory[16'h7ed6] <= 8'h5c;
		memory[16'h7ed7] <= 8'h77;
		memory[16'h7ed8] <= 8'hcc;
		memory[16'h7ed9] <= 8'ha2;
		memory[16'h7eda] <= 8'h5f;
		memory[16'h7edb] <= 8'h45;
		memory[16'h7edc] <= 8'hf0;
		memory[16'h7edd] <= 8'h95;
		memory[16'h7ede] <= 8'h86;
		memory[16'h7edf] <= 8'h82;
		memory[16'h7ee0] <= 8'h58;
		memory[16'h7ee1] <= 8'hc0;
		memory[16'h7ee2] <= 8'h45;
		memory[16'h7ee3] <= 8'had;
		memory[16'h7ee4] <= 8'h8e;
		memory[16'h7ee5] <= 8'h0;
		memory[16'h7ee6] <= 8'hbd;
		memory[16'h7ee7] <= 8'h48;
		memory[16'h7ee8] <= 8'hd3;
		memory[16'h7ee9] <= 8'hfd;
		memory[16'h7eea] <= 8'h5c;
		memory[16'h7eeb] <= 8'h17;
		memory[16'h7eec] <= 8'hfe;
		memory[16'h7eed] <= 8'h41;
		memory[16'h7eee] <= 8'h77;
		memory[16'h7eef] <= 8'hcb;
		memory[16'h7ef0] <= 8'h1b;
		memory[16'h7ef1] <= 8'h8;
		memory[16'h7ef2] <= 8'h6f;
		memory[16'h7ef3] <= 8'hb9;
		memory[16'h7ef4] <= 8'h94;
		memory[16'h7ef5] <= 8'hcb;
		memory[16'h7ef6] <= 8'h30;
		memory[16'h7ef7] <= 8'h61;
		memory[16'h7ef8] <= 8'h6d;
		memory[16'h7ef9] <= 8'h90;
		memory[16'h7efa] <= 8'ha6;
		memory[16'h7efb] <= 8'h5e;
		memory[16'h7efc] <= 8'h25;
		memory[16'h7efd] <= 8'h2c;
		memory[16'h7efe] <= 8'he0;
		memory[16'h7eff] <= 8'h7d;
		memory[16'h7f00] <= 8'hed;
		memory[16'h7f01] <= 8'h25;
		memory[16'h7f02] <= 8'h2a;
		memory[16'h7f03] <= 8'h7b;
		memory[16'h7f04] <= 8'h26;
		memory[16'h7f05] <= 8'he8;
		memory[16'h7f06] <= 8'hc3;
		memory[16'h7f07] <= 8'hf9;
		memory[16'h7f08] <= 8'he5;
		memory[16'h7f09] <= 8'h20;
		memory[16'h7f0a] <= 8'h11;
		memory[16'h7f0b] <= 8'he3;
		memory[16'h7f0c] <= 8'h61;
		memory[16'h7f0d] <= 8'h88;
		memory[16'h7f0e] <= 8'haf;
		memory[16'h7f0f] <= 8'h7c;
		memory[16'h7f10] <= 8'h90;
		memory[16'h7f11] <= 8'h1e;
		memory[16'h7f12] <= 8'h35;
		memory[16'h7f13] <= 8'h25;
		memory[16'h7f14] <= 8'he9;
		memory[16'h7f15] <= 8'h66;
		memory[16'h7f16] <= 8'h86;
		memory[16'h7f17] <= 8'h57;
		memory[16'h7f18] <= 8'hf6;
		memory[16'h7f19] <= 8'h2c;
		memory[16'h7f1a] <= 8'hb5;
		memory[16'h7f1b] <= 8'h1b;
		memory[16'h7f1c] <= 8'h59;
		memory[16'h7f1d] <= 8'h95;
		memory[16'h7f1e] <= 8'h98;
		memory[16'h7f1f] <= 8'h46;
		memory[16'h7f20] <= 8'hbb;
		memory[16'h7f21] <= 8'hc2;
		memory[16'h7f22] <= 8'hc1;
		memory[16'h7f23] <= 8'he1;
		memory[16'h7f24] <= 8'haa;
		memory[16'h7f25] <= 8'h85;
		memory[16'h7f26] <= 8'hda;
		memory[16'h7f27] <= 8'h90;
		memory[16'h7f28] <= 8'ha5;
		memory[16'h7f29] <= 8'heb;
		memory[16'h7f2a] <= 8'h73;
		memory[16'h7f2b] <= 8'h6;
		memory[16'h7f2c] <= 8'h74;
		memory[16'h7f2d] <= 8'h22;
		memory[16'h7f2e] <= 8'h83;
		memory[16'h7f2f] <= 8'h4;
		memory[16'h7f30] <= 8'h40;
		memory[16'h7f31] <= 8'hb8;
		memory[16'h7f32] <= 8'h29;
		memory[16'h7f33] <= 8'h2a;
		memory[16'h7f34] <= 8'h1e;
		memory[16'h7f35] <= 8'haf;
		memory[16'h7f36] <= 8'h81;
		memory[16'h7f37] <= 8'h14;
		memory[16'h7f38] <= 8'hdc;
		memory[16'h7f39] <= 8'h36;
		memory[16'h7f3a] <= 8'h2f;
		memory[16'h7f3b] <= 8'h35;
		memory[16'h7f3c] <= 8'hcb;
		memory[16'h7f3d] <= 8'hc7;
		memory[16'h7f3e] <= 8'h7b;
		memory[16'h7f3f] <= 8'h86;
		memory[16'h7f40] <= 8'h8a;
		memory[16'h7f41] <= 8'h3c;
		memory[16'h7f42] <= 8'h67;
		memory[16'h7f43] <= 8'h34;
		memory[16'h7f44] <= 8'hc1;
		memory[16'h7f45] <= 8'h42;
		memory[16'h7f46] <= 8'hc4;
		memory[16'h7f47] <= 8'h66;
		memory[16'h7f48] <= 8'h2d;
		memory[16'h7f49] <= 8'h38;
		memory[16'h7f4a] <= 8'h6d;
		memory[16'h7f4b] <= 8'ha1;
		memory[16'h7f4c] <= 8'h5a;
		memory[16'h7f4d] <= 8'hf0;
		memory[16'h7f4e] <= 8'ha6;
		memory[16'h7f4f] <= 8'h9b;
		memory[16'h7f50] <= 8'ha8;
		memory[16'h7f51] <= 8'hcf;
		memory[16'h7f52] <= 8'hc5;
		memory[16'h7f53] <= 8'hc7;
		memory[16'h7f54] <= 8'h7f;
		memory[16'h7f55] <= 8'h46;
		memory[16'h7f56] <= 8'hdb;
		memory[16'h7f57] <= 8'h5b;
		memory[16'h7f58] <= 8'h7c;
		memory[16'h7f59] <= 8'hb;
		memory[16'h7f5a] <= 8'h90;
		memory[16'h7f5b] <= 8'h47;
		memory[16'h7f5c] <= 8'hd2;
		memory[16'h7f5d] <= 8'hb;
		memory[16'h7f5e] <= 8'hce;
		memory[16'h7f5f] <= 8'h5c;
		memory[16'h7f60] <= 8'h47;
		memory[16'h7f61] <= 8'h35;
		memory[16'h7f62] <= 8'h91;
		memory[16'h7f63] <= 8'h9;
		memory[16'h7f64] <= 8'h77;
		memory[16'h7f65] <= 8'h55;
		memory[16'h7f66] <= 8'h6f;
		memory[16'h7f67] <= 8'ha5;
		memory[16'h7f68] <= 8'h8d;
		memory[16'h7f69] <= 8'hdc;
		memory[16'h7f6a] <= 8'h46;
		memory[16'h7f6b] <= 8'he8;
		memory[16'h7f6c] <= 8'hcc;
		memory[16'h7f6d] <= 8'hec;
		memory[16'h7f6e] <= 8'h83;
		memory[16'h7f6f] <= 8'h75;
		memory[16'h7f70] <= 8'hbc;
		memory[16'h7f71] <= 8'h48;
		memory[16'h7f72] <= 8'h3c;
		memory[16'h7f73] <= 8'h3b;
		memory[16'h7f74] <= 8'h8e;
		memory[16'h7f75] <= 8'h17;
		memory[16'h7f76] <= 8'h96;
		memory[16'h7f77] <= 8'ha;
		memory[16'h7f78] <= 8'h22;
		memory[16'h7f79] <= 8'h26;
		memory[16'h7f7a] <= 8'h51;
		memory[16'h7f7b] <= 8'hf5;
		memory[16'h7f7c] <= 8'h31;
		memory[16'h7f7d] <= 8'h1f;
		memory[16'h7f7e] <= 8'h51;
		memory[16'h7f7f] <= 8'h78;
		memory[16'h7f80] <= 8'h55;
		memory[16'h7f81] <= 8'he2;
		memory[16'h7f82] <= 8'h81;
		memory[16'h7f83] <= 8'hcc;
		memory[16'h7f84] <= 8'h38;
		memory[16'h7f85] <= 8'hf1;
		memory[16'h7f86] <= 8'h71;
		memory[16'h7f87] <= 8'hc5;
		memory[16'h7f88] <= 8'hcd;
		memory[16'h7f89] <= 8'hb8;
		memory[16'h7f8a] <= 8'had;
		memory[16'h7f8b] <= 8'h9a;
		memory[16'h7f8c] <= 8'ha4;
		memory[16'h7f8d] <= 8'h30;
		memory[16'h7f8e] <= 8'hf;
		memory[16'h7f8f] <= 8'h60;
		memory[16'h7f90] <= 8'h78;
		memory[16'h7f91] <= 8'h4b;
		memory[16'h7f92] <= 8'h9b;
		memory[16'h7f93] <= 8'h6;
		memory[16'h7f94] <= 8'h62;
		memory[16'h7f95] <= 8'h31;
		memory[16'h7f96] <= 8'h10;
		memory[16'h7f97] <= 8'h85;
		memory[16'h7f98] <= 8'h57;
		memory[16'h7f99] <= 8'h62;
		memory[16'h7f9a] <= 8'h7a;
		memory[16'h7f9b] <= 8'h88;
		memory[16'h7f9c] <= 8'h81;
		memory[16'h7f9d] <= 8'hcb;
		memory[16'h7f9e] <= 8'h1;
		memory[16'h7f9f] <= 8'hd6;
		memory[16'h7fa0] <= 8'hae;
		memory[16'h7fa1] <= 8'h82;
		memory[16'h7fa2] <= 8'ha3;
		memory[16'h7fa3] <= 8'he6;
		memory[16'h7fa4] <= 8'h73;
		memory[16'h7fa5] <= 8'h14;
		memory[16'h7fa6] <= 8'hab;
		memory[16'h7fa7] <= 8'h41;
		memory[16'h7fa8] <= 8'hcc;
		memory[16'h7fa9] <= 8'h59;
		memory[16'h7faa] <= 8'hdb;
		memory[16'h7fab] <= 8'h71;
		memory[16'h7fac] <= 8'h89;
		memory[16'h7fad] <= 8'hea;
		memory[16'h7fae] <= 8'hd1;
		memory[16'h7faf] <= 8'h2;
		memory[16'h7fb0] <= 8'h35;
		memory[16'h7fb1] <= 8'h6d;
		memory[16'h7fb2] <= 8'h8;
		memory[16'h7fb3] <= 8'h97;
		memory[16'h7fb4] <= 8'h9e;
		memory[16'h7fb5] <= 8'h19;
		memory[16'h7fb6] <= 8'h1c;
		memory[16'h7fb7] <= 8'hf6;
		memory[16'h7fb8] <= 8'h7b;
		memory[16'h7fb9] <= 8'h96;
		memory[16'h7fba] <= 8'h7e;
		memory[16'h7fbb] <= 8'hfc;
		memory[16'h7fbc] <= 8'h62;
		memory[16'h7fbd] <= 8'h7f;
		memory[16'h7fbe] <= 8'hd3;
		memory[16'h7fbf] <= 8'h10;
		memory[16'h7fc0] <= 8'h2;
		memory[16'h7fc1] <= 8'h76;
		memory[16'h7fc2] <= 8'hf6;
		memory[16'h7fc3] <= 8'h75;
		memory[16'h7fc4] <= 8'h8a;
		memory[16'h7fc5] <= 8'ha1;
		memory[16'h7fc6] <= 8'hb6;
		memory[16'h7fc7] <= 8'h57;
		memory[16'h7fc8] <= 8'hfa;
		memory[16'h7fc9] <= 8'h91;
		memory[16'h7fca] <= 8'hc8;
		memory[16'h7fcb] <= 8'h84;
		memory[16'h7fcc] <= 8'h7b;
		memory[16'h7fcd] <= 8'h99;
		memory[16'h7fce] <= 8'h86;
		memory[16'h7fcf] <= 8'hb0;
		memory[16'h7fd0] <= 8'h6;
		memory[16'h7fd1] <= 8'h8e;
		memory[16'h7fd2] <= 8'h48;
		memory[16'h7fd3] <= 8'ha5;
		memory[16'h7fd4] <= 8'ha7;
		memory[16'h7fd5] <= 8'h64;
		memory[16'h7fd6] <= 8'h9b;
		memory[16'h7fd7] <= 8'h22;
		memory[16'h7fd8] <= 8'hfb;
		memory[16'h7fd9] <= 8'h19;
		memory[16'h7fda] <= 8'h1f;
		memory[16'h7fdb] <= 8'h5d;
		memory[16'h7fdc] <= 8'h99;
		memory[16'h7fdd] <= 8'hf2;
		memory[16'h7fde] <= 8'h6d;
		memory[16'h7fdf] <= 8'h9b;
		memory[16'h7fe0] <= 8'h68;
		memory[16'h7fe1] <= 8'h63;
		memory[16'h7fe2] <= 8'h10;
		memory[16'h7fe3] <= 8'hf2;
		memory[16'h7fe4] <= 8'h4;
		memory[16'h7fe5] <= 8'hc7;
		memory[16'h7fe6] <= 8'h49;
		memory[16'h7fe7] <= 8'hff;
		memory[16'h7fe8] <= 8'h58;
		memory[16'h7fe9] <= 8'h11;
		memory[16'h7fea] <= 8'h83;
		memory[16'h7feb] <= 8'hd4;
		memory[16'h7fec] <= 8'hab;
		memory[16'h7fed] <= 8'h9;
		memory[16'h7fee] <= 8'h84;
		memory[16'h7fef] <= 8'hb1;
		memory[16'h7ff0] <= 8'h97;
		memory[16'h7ff1] <= 8'hcc;
		memory[16'h7ff2] <= 8'h56;
		memory[16'h7ff3] <= 8'h3f;
		memory[16'h7ff4] <= 8'h31;
		memory[16'h7ff5] <= 8'hf1;
		memory[16'h7ff6] <= 8'h61;
		memory[16'h7ff7] <= 8'h2c;
		memory[16'h7ff8] <= 8'hb;
		memory[16'h7ff9] <= 8'h80;
		memory[16'h7ffa] <= 8'h89;
		memory[16'h7ffb] <= 8'ha4;
		memory[16'h7ffc] <= 8'h72;
		memory[16'h7ffd] <= 8'hf6;
		memory[16'h7ffe] <= 8'h3f;
		memory[16'h7fff] <= 8'hda;
	end
endmodule
