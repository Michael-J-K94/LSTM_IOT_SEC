`timescale 1ns/100ps
`define INIT_DELAY 10
`define INTERVAL 1
`define MEM_SIZE 65536

module br_bias_memory(
	input readM,
	output reg ready,
	output reg [7:0] data
	);

	reg [7:0] memory [`MEM_SIZE - 1:0];
	reg [15:0] address;

	always begin
		#`INIT_DELAY
		forever begin
			wait(readM == 1);
			#`INTERVAL;
			data = memory[address];
			address = address + 1;
			ready = 1;
			wait(readM == 0);
			#`INTERVAL;
			ready = 0;
		end
	end

	initial begin
		address <= 0;
		ready <= 0;
	end

	initial begin
		memory[16'h0] <= 8'h80;
		memory[16'h1] <= 8'h80;
		memory[16'h2] <= 8'h80;
		memory[16'h3] <= 8'h80;
		memory[16'h4] <= 8'h80;
		memory[16'h5] <= 8'h80;
		memory[16'h6] <= 8'h80;
		memory[16'h7] <= 8'h80;
		memory[16'h8] <= 8'h80;
		memory[16'h9] <= 8'h80;
		memory[16'ha] <= 8'h80;
		memory[16'hb] <= 8'h80;
		memory[16'hc] <= 8'h80;
		memory[16'hd] <= 8'h80;
		memory[16'he] <= 8'h80;
		memory[16'hf] <= 8'h80;
		memory[16'h10] <= 8'h80;
		memory[16'h11] <= 8'h80;
		memory[16'h12] <= 8'h80;
		memory[16'h13] <= 8'h80;
		memory[16'h14] <= 8'h80;
		memory[16'h15] <= 8'h80;
		memory[16'h16] <= 8'h80;
		memory[16'h17] <= 8'h80;
		memory[16'h18] <= 8'h80;
		memory[16'h19] <= 8'h80;
		memory[16'h1a] <= 8'h80;
		memory[16'h1b] <= 8'h80;
		memory[16'h1c] <= 8'h80;
		memory[16'h1d] <= 8'h80;
		memory[16'h1e] <= 8'h80;
		memory[16'h1f] <= 8'h80;
		memory[16'h20] <= 8'h80;
		memory[16'h21] <= 8'h80;
		memory[16'h22] <= 8'h80;
		memory[16'h23] <= 8'h80;
		memory[16'h24] <= 8'h80;
		memory[16'h25] <= 8'h80;
		memory[16'h26] <= 8'h80;
		memory[16'h27] <= 8'h80;
		memory[16'h28] <= 8'h80;
		memory[16'h29] <= 8'h80;
		memory[16'h2a] <= 8'h80;
		memory[16'h2b] <= 8'h80;
		memory[16'h2c] <= 8'h80;
		memory[16'h2d] <= 8'h80;
		memory[16'h2e] <= 8'h80;
		memory[16'h2f] <= 8'h80;
		memory[16'h30] <= 8'h80;
		memory[16'h31] <= 8'h80;
		memory[16'h32] <= 8'h80;
		memory[16'h33] <= 8'h80;
		memory[16'h34] <= 8'h80;
		memory[16'h35] <= 8'h80;
		memory[16'h36] <= 8'h80;
		memory[16'h37] <= 8'h80;
		memory[16'h38] <= 8'h80;
		memory[16'h39] <= 8'h80;
		memory[16'h3a] <= 8'h80;
		memory[16'h3b] <= 8'h80;
		memory[16'h3c] <= 8'h80;
		memory[16'h3d] <= 8'h80;
		memory[16'h3e] <= 8'h80;
		memory[16'h3f] <= 8'h80;
		memory[16'h40] <= 8'h80;
		memory[16'h41] <= 8'h80;
		memory[16'h42] <= 8'h80;
		memory[16'h43] <= 8'h80;
		memory[16'h44] <= 8'h80;
		memory[16'h45] <= 8'h80;
		memory[16'h46] <= 8'h80;
		memory[16'h47] <= 8'h80;
		memory[16'h48] <= 8'h80;
		memory[16'h49] <= 8'h80;
		memory[16'h4a] <= 8'h80;
		memory[16'h4b] <= 8'h80;
		memory[16'h4c] <= 8'h80;
		memory[16'h4d] <= 8'h80;
		memory[16'h4e] <= 8'h80;
		memory[16'h4f] <= 8'h80;
		memory[16'h50] <= 8'h80;
		memory[16'h51] <= 8'h80;
		memory[16'h52] <= 8'h80;
		memory[16'h53] <= 8'h80;
		memory[16'h54] <= 8'h80;
		memory[16'h55] <= 8'h80;
		memory[16'h56] <= 8'h80;
		memory[16'h57] <= 8'h80;
		memory[16'h58] <= 8'h80;
		memory[16'h59] <= 8'h80;
		memory[16'h5a] <= 8'h80;
		memory[16'h5b] <= 8'h80;
		memory[16'h5c] <= 8'h80;
		memory[16'h5d] <= 8'h80;
		memory[16'h5e] <= 8'h80;
		memory[16'h5f] <= 8'h80;
		memory[16'h60] <= 8'h80;
		memory[16'h61] <= 8'h80;
		memory[16'h62] <= 8'h80;
		memory[16'h63] <= 8'h80;
		memory[16'h64] <= 8'h80;
		memory[16'h65] <= 8'h80;
		memory[16'h66] <= 8'h80;
		memory[16'h67] <= 8'h80;
		memory[16'h68] <= 8'h80;
		memory[16'h69] <= 8'h80;
		memory[16'h6a] <= 8'h80;
		memory[16'h6b] <= 8'h80;
		memory[16'h6c] <= 8'h80;
		memory[16'h6d] <= 8'h80;
		memory[16'h6e] <= 8'h80;
		memory[16'h6f] <= 8'h80;
		memory[16'h70] <= 8'h80;
		memory[16'h71] <= 8'h80;
		memory[16'h72] <= 8'h80;
		memory[16'h73] <= 8'h80;
		memory[16'h74] <= 8'h80;
		memory[16'h75] <= 8'h80;
		memory[16'h76] <= 8'h80;
		memory[16'h77] <= 8'h80;
		memory[16'h78] <= 8'h80;
		memory[16'h79] <= 8'h80;
		memory[16'h7a] <= 8'h80;
		memory[16'h7b] <= 8'h80;
		memory[16'h7c] <= 8'h80;
		memory[16'h7d] <= 8'h80;
		memory[16'h7e] <= 8'h80;
		memory[16'h7f] <= 8'h80;
		memory[16'h80] <= 8'h80;
		memory[16'h81] <= 8'h80;
		memory[16'h82] <= 8'h80;
		memory[16'h83] <= 8'h80;
		memory[16'h84] <= 8'h80;
		memory[16'h85] <= 8'h80;
		memory[16'h86] <= 8'h80;
		memory[16'h87] <= 8'h80;
		memory[16'h88] <= 8'h80;
		memory[16'h89] <= 8'h80;
		memory[16'h8a] <= 8'h80;
		memory[16'h8b] <= 8'h80;
		memory[16'h8c] <= 8'h80;
		memory[16'h8d] <= 8'h80;
		memory[16'h8e] <= 8'h80;
		memory[16'h8f] <= 8'h80;
		memory[16'h90] <= 8'h80;
		memory[16'h91] <= 8'h80;
		memory[16'h92] <= 8'h80;
		memory[16'h93] <= 8'h80;
		memory[16'h94] <= 8'h80;
		memory[16'h95] <= 8'h80;
		memory[16'h96] <= 8'h80;
		memory[16'h97] <= 8'h80;
		memory[16'h98] <= 8'h80;
		memory[16'h99] <= 8'h80;
		memory[16'h9a] <= 8'h80;
		memory[16'h9b] <= 8'h80;
		memory[16'h9c] <= 8'h80;
		memory[16'h9d] <= 8'h80;
		memory[16'h9e] <= 8'h80;
		memory[16'h9f] <= 8'h80;
		memory[16'ha0] <= 8'h80;
		memory[16'ha1] <= 8'h80;
		memory[16'ha2] <= 8'h80;
		memory[16'ha3] <= 8'h80;
		memory[16'ha4] <= 8'h80;
		memory[16'ha5] <= 8'h80;
		memory[16'ha6] <= 8'h80;
		memory[16'ha7] <= 8'h80;
		memory[16'ha8] <= 8'h80;
		memory[16'ha9] <= 8'h80;
		memory[16'haa] <= 8'h80;
		memory[16'hab] <= 8'h80;
		memory[16'hac] <= 8'h80;
		memory[16'had] <= 8'h80;
		memory[16'hae] <= 8'h80;
		memory[16'haf] <= 8'h80;
		memory[16'hb0] <= 8'h80;
		memory[16'hb1] <= 8'h80;
		memory[16'hb2] <= 8'h80;
		memory[16'hb3] <= 8'h80;
		memory[16'hb4] <= 8'h80;
		memory[16'hb5] <= 8'h80;
		memory[16'hb6] <= 8'h80;
		memory[16'hb7] <= 8'h80;
		memory[16'hb8] <= 8'h80;
		memory[16'hb9] <= 8'h80;
		memory[16'hba] <= 8'h80;
		memory[16'hbb] <= 8'h80;
		memory[16'hbc] <= 8'h80;
		memory[16'hbd] <= 8'h80;
		memory[16'hbe] <= 8'h80;
		memory[16'hbf] <= 8'h80;
		memory[16'hc0] <= 8'h80;
		memory[16'hc1] <= 8'h80;
		memory[16'hc2] <= 8'h80;
		memory[16'hc3] <= 8'h80;
		memory[16'hc4] <= 8'h80;
		memory[16'hc5] <= 8'h80;
		memory[16'hc6] <= 8'h80;
		memory[16'hc7] <= 8'h80;
		memory[16'hc8] <= 8'h80;
		memory[16'hc9] <= 8'h80;
		memory[16'hca] <= 8'h80;
		memory[16'hcb] <= 8'h80;
		memory[16'hcc] <= 8'h80;
		memory[16'hcd] <= 8'h80;
		memory[16'hce] <= 8'h80;
		memory[16'hcf] <= 8'h80;
		memory[16'hd0] <= 8'h80;
		memory[16'hd1] <= 8'h80;
		memory[16'hd2] <= 8'h80;
		memory[16'hd3] <= 8'h80;
		memory[16'hd4] <= 8'h80;
		memory[16'hd5] <= 8'h80;
		memory[16'hd6] <= 8'h80;
		memory[16'hd7] <= 8'h80;
		memory[16'hd8] <= 8'h80;
		memory[16'hd9] <= 8'h80;
		memory[16'hda] <= 8'h80;
		memory[16'hdb] <= 8'h80;
		memory[16'hdc] <= 8'h80;
		memory[16'hdd] <= 8'h80;
		memory[16'hde] <= 8'h80;
		memory[16'hdf] <= 8'h80;
		memory[16'he0] <= 8'h80;
		memory[16'he1] <= 8'h80;
		memory[16'he2] <= 8'h80;
		memory[16'he3] <= 8'h80;
		memory[16'he4] <= 8'h80;
		memory[16'he5] <= 8'h80;
		memory[16'he6] <= 8'h80;
		memory[16'he7] <= 8'h80;
		memory[16'he8] <= 8'h80;
		memory[16'he9] <= 8'h80;
		memory[16'hea] <= 8'h80;
		memory[16'heb] <= 8'h80;
		memory[16'hec] <= 8'h80;
		memory[16'hed] <= 8'h80;
		memory[16'hee] <= 8'h80;
		memory[16'hef] <= 8'h80;
		memory[16'hf0] <= 8'h80;
		memory[16'hf1] <= 8'h80;
		memory[16'hf2] <= 8'h80;
		memory[16'hf3] <= 8'h80;
		memory[16'hf4] <= 8'h80;
		memory[16'hf5] <= 8'h80;
		memory[16'hf6] <= 8'h80;
		memory[16'hf7] <= 8'h80;
		memory[16'hf8] <= 8'h80;
		memory[16'hf9] <= 8'h80;
		memory[16'hfa] <= 8'h80;
		memory[16'hfb] <= 8'h80;
		memory[16'hfc] <= 8'h80;
		memory[16'hfd] <= 8'h80;
		memory[16'hfe] <= 8'h80;
		memory[16'hff] <= 8'h80;
	end
endmodule
